-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant foo_base_address : std_logic_vector(3 downto 0) := "0000";
  constant free_queue_base_address : std_logic_vector(2 downto 0) := "000";
  constant free_queue_ram_base_address : std_logic_vector(10 downto 0) := "00000000001";
  constant mempool_base_address : std_logic_vector(10 downto 0) := "00000000000";
  constant xx_xstr1_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr2_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr3_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr4_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr5_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr6_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr7_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr8_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr_base_address : std_logic_vector(4 downto 0) := "00000";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_foo is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_foo;
architecture Default of default_initializer_foo is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_foo_CP_217_start: Boolean;
  -- links between control-path and data-path
  signal binary_156_inst_req_0 : boolean;
  signal binary_156_inst_ack_0 : boolean;
  signal binary_156_inst_req_1 : boolean;
  signal binary_156_inst_ack_1 : boolean;
  signal array_obj_ref_159_index_0_resize_req_0 : boolean;
  signal array_obj_ref_159_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_159_index_0_rename_req_0 : boolean;
  signal array_obj_ref_159_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_159_offset_inst_req_0 : boolean;
  signal array_obj_ref_159_offset_inst_ack_0 : boolean;
  signal array_obj_ref_159_root_address_inst_req_0 : boolean;
  signal array_obj_ref_159_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_159_addr_0_req_0 : boolean;
  signal array_obj_ref_159_addr_0_ack_0 : boolean;
  signal array_obj_ref_159_gather_scatter_req_0 : boolean;
  signal array_obj_ref_159_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_159_store_0_req_0 : boolean;
  signal array_obj_ref_159_store_0_ack_0 : boolean;
  signal array_obj_ref_159_store_0_req_1 : boolean;
  signal array_obj_ref_159_store_0_ack_1 : boolean;
  signal binary_165_inst_req_0 : boolean;
  signal binary_165_inst_ack_0 : boolean;
  signal binary_165_inst_req_1 : boolean;
  signal binary_165_inst_ack_1 : boolean;
  signal if_stmt_162_branch_req_0 : boolean;
  signal if_stmt_162_branch_ack_1 : boolean;
  signal if_stmt_162_branch_ack_0 : boolean;
  signal phi_stmt_146_req_0 : boolean;
  signal phi_stmt_146_req_1 : boolean;
  signal phi_stmt_146_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_foo_CP_217: Block -- control-path 
    signal cp_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(30) & cp_elements(26));
    binary_156_inst_req_0 <= cp_elements(1);
    cp_elements(2) <= OrReduce(cp_elements(15) & cp_elements(23));
    cp_elements(3) <= binary_156_inst_ack_0;
    binary_156_inst_req_1 <= cp_elements(3);
    cp_elements(4) <= binary_156_inst_ack_1;
    array_obj_ref_159_index_0_resize_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_159_index_0_resize_ack_0;
    array_obj_ref_159_index_0_rename_req_0 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_159_index_0_rename_ack_0;
    array_obj_ref_159_offset_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_159_offset_inst_ack_0;
    array_obj_ref_159_root_address_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_159_root_address_inst_ack_0;
    array_obj_ref_159_addr_0_req_0 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_159_addr_0_ack_0;
    array_obj_ref_159_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_159_gather_scatter_ack_0;
    array_obj_ref_159_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_159_store_0_ack_0;
    array_obj_ref_159_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_159_store_0_ack_1;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= false;
    cp_elements(15) <= cp_elements(14);
    cp_elements(16) <= cp_elements(12);
    binary_165_inst_req_0 <= cp_elements(16);
    cp_elements(17) <= binary_165_inst_ack_0;
    binary_165_inst_req_1 <= cp_elements(17);
    cp_elements(18) <= binary_165_inst_ack_1;
    if_stmt_162_branch_req_0 <= cp_elements(18);
    cp_elements(19) <= cp_elements(18);
    cp_elements(20) <= cp_elements(19);
    cp_elements(21) <= if_stmt_162_branch_ack_1;
    phi_stmt_146_req_1 <= cp_elements(21);
    cp_elements(22) <= cp_elements(19);
    cp_elements(23) <= if_stmt_162_branch_ack_0;
    cp_elements(24) <= cp_elements(0);
    cp_elements(25) <= false;
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(0);
    phi_stmt_146_req_0 <= cp_elements(27);
    cp_elements(28) <= OrReduce(cp_elements(27) & cp_elements(21));
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= phi_stmt_146_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_0_146 : std_logic_vector(3 downto 0);
    signal array_obj_ref_159_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_159_final_offset : std_logic_vector(3 downto 0);
    signal array_obj_ref_159_offset_scale_factor_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_159_resized_base_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_159_root_address : std_logic_vector(3 downto 0);
    signal array_obj_ref_159_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_159_word_offset_0 : std_logic_vector(3 downto 0);
    signal binary_165_wire : std_logic_vector(0 downto 0);
    signal expr_155_wire_constant : std_logic_vector(3 downto 0);
    signal expr_160_wire_constant : std_logic_vector(7 downto 0);
    signal expr_164_wire_constant : std_logic_vector(3 downto 0);
    signal next_I_157 : std_logic_vector(3 downto 0);
    signal simple_obj_ref_158_resized : std_logic_vector(3 downto 0);
    signal simple_obj_ref_158_scaled : std_logic_vector(3 downto 0);
    signal type_cast_150_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    array_obj_ref_159_offset_scale_factor_0 <= "0001";
    array_obj_ref_159_resized_base_address <= "0000";
    array_obj_ref_159_word_offset_0 <= "0000";
    expr_155_wire_constant <= "0001";
    expr_160_wire_constant <= "00000000";
    expr_164_wire_constant <= "1010";
    type_cast_150_wire_constant <= "0000";
    phi_stmt_146: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_150_wire_constant & next_I_157;
      req <= phi_stmt_146_req_0 & phi_stmt_146_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_146_ack_0,
          idata => idata,
          odata => I_0_146,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_146
    array_obj_ref_159_index_0_resize: RegisterBase --
      generic map(in_data_width => 4,out_data_width => 4, flow_through => true ) 
      port map( din => I_0_146, dout => simple_obj_ref_158_resized, req => array_obj_ref_159_index_0_resize_req_0, ack => array_obj_ref_159_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_159_offset_inst: RegisterBase --
      generic map(in_data_width => 4,out_data_width => 4, flow_through => true ) 
      port map( din => simple_obj_ref_158_scaled, dout => array_obj_ref_159_final_offset, req => array_obj_ref_159_offset_inst_req_0, ack => array_obj_ref_159_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_159_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(3 downto 0); --
    begin -- 
      array_obj_ref_159_addr_0_ack_0 <= array_obj_ref_159_addr_0_req_0;
      aggregated_sig <= array_obj_ref_159_root_address;
      array_obj_ref_159_word_address_0 <= aggregated_sig(3 downto 0);
      --
    end Block;
    array_obj_ref_159_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_159_gather_scatter_ack_0 <= array_obj_ref_159_gather_scatter_req_0;
      aggregated_sig <= expr_160_wire_constant;
      array_obj_ref_159_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_159_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(3 downto 0); --
    begin -- 
      array_obj_ref_159_index_0_rename_ack_0 <= array_obj_ref_159_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_158_resized;
      simple_obj_ref_158_scaled <= aggregated_sig(3 downto 0);
      --
    end Block;
    array_obj_ref_159_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(3 downto 0); --
    begin -- 
      array_obj_ref_159_root_address_inst_ack_0 <= array_obj_ref_159_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_159_final_offset;
      array_obj_ref_159_root_address <= aggregated_sig(3 downto 0);
      --
    end Block;
    if_stmt_162_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_165_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_162_branch_req_0,
          ack0 => if_stmt_162_branch_ack_0,
          ack1 => if_stmt_162_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_156_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(3 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_0_146;
      next_I_157 <= data_out(3 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 4,
          constant_operand => "0001",
          constant_width => 4,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_156_inst_req_0,
          ackL => binary_156_inst_ack_0,
          reqR => binary_156_inst_req_1,
          ackR => binary_156_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_165_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= next_I_157;
      binary_165_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 4,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "1010",
          constant_width => 4,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_165_inst_req_0,
          ackL => binary_165_inst_ack_0,
          reqR => binary_165_inst_req_1,
          ackR => binary_165_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_159_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_159_store_0_req_0;
      array_obj_ref_159_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_159_store_0_req_1;
      array_obj_ref_159_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_159_word_address_0;
      data_in <= array_obj_ref_159_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(3 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_free_queue is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_free_queue;
architecture Default of default_initializer_free_queue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_free_queue_CP_351_start: Boolean;
  -- links between control-path and data-path
  signal binary_185_inst_req_0 : boolean;
  signal binary_185_inst_ack_0 : boolean;
  signal binary_185_inst_req_1 : boolean;
  signal binary_185_inst_ack_1 : boolean;
  signal array_obj_ref_188_index_0_resize_req_0 : boolean;
  signal array_obj_ref_188_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_188_index_0_rename_req_0 : boolean;
  signal array_obj_ref_188_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_188_offset_inst_req_0 : boolean;
  signal array_obj_ref_188_offset_inst_ack_0 : boolean;
  signal array_obj_ref_188_root_address_inst_req_0 : boolean;
  signal array_obj_ref_188_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_188_addr_0_req_0 : boolean;
  signal array_obj_ref_188_addr_0_ack_0 : boolean;
  signal array_obj_ref_188_gather_scatter_req_0 : boolean;
  signal array_obj_ref_188_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_188_store_0_req_0 : boolean;
  signal array_obj_ref_188_store_0_ack_0 : boolean;
  signal array_obj_ref_188_store_0_req_1 : boolean;
  signal array_obj_ref_188_store_0_ack_1 : boolean;
  signal binary_194_inst_req_0 : boolean;
  signal binary_194_inst_ack_0 : boolean;
  signal binary_194_inst_req_1 : boolean;
  signal binary_194_inst_ack_1 : boolean;
  signal if_stmt_191_branch_req_0 : boolean;
  signal if_stmt_191_branch_ack_1 : boolean;
  signal if_stmt_191_branch_ack_0 : boolean;
  signal phi_stmt_175_req_0 : boolean;
  signal phi_stmt_175_req_1 : boolean;
  signal phi_stmt_175_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_free_queue_CP_351: Block -- control-path 
    signal cp_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(26) & cp_elements(30));
    binary_185_inst_req_0 <= cp_elements(1);
    cp_elements(2) <= OrReduce(cp_elements(23) & cp_elements(15));
    cp_elements(3) <= binary_185_inst_ack_0;
    binary_185_inst_req_1 <= cp_elements(3);
    cp_elements(4) <= binary_185_inst_ack_1;
    array_obj_ref_188_index_0_resize_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_188_index_0_resize_ack_0;
    array_obj_ref_188_index_0_rename_req_0 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_188_index_0_rename_ack_0;
    array_obj_ref_188_offset_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_188_offset_inst_ack_0;
    array_obj_ref_188_root_address_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_188_root_address_inst_ack_0;
    array_obj_ref_188_addr_0_req_0 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_188_addr_0_ack_0;
    array_obj_ref_188_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_188_gather_scatter_ack_0;
    array_obj_ref_188_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_188_store_0_ack_0;
    array_obj_ref_188_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_188_store_0_ack_1;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= false;
    cp_elements(15) <= cp_elements(14);
    cp_elements(16) <= cp_elements(12);
    binary_194_inst_req_0 <= cp_elements(16);
    cp_elements(17) <= binary_194_inst_ack_0;
    binary_194_inst_req_1 <= cp_elements(17);
    cp_elements(18) <= binary_194_inst_ack_1;
    if_stmt_191_branch_req_0 <= cp_elements(18);
    cp_elements(19) <= cp_elements(18);
    cp_elements(20) <= cp_elements(19);
    cp_elements(21) <= if_stmt_191_branch_ack_1;
    phi_stmt_175_req_1 <= cp_elements(21);
    cp_elements(22) <= cp_elements(19);
    cp_elements(23) <= if_stmt_191_branch_ack_0;
    cp_elements(24) <= cp_elements(0);
    cp_elements(25) <= false;
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(0);
    phi_stmt_175_req_0 <= cp_elements(27);
    cp_elements(28) <= OrReduce(cp_elements(21) & cp_elements(27));
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= phi_stmt_175_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_0_175 : std_logic_vector(2 downto 0);
    signal array_obj_ref_188_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_188_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_188_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_188_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_188_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_188_word_address_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_188_word_offset_0 : std_logic_vector(2 downto 0);
    signal binary_194_wire : std_logic_vector(0 downto 0);
    signal expr_184_wire_constant : std_logic_vector(2 downto 0);
    signal expr_189_wire_constant : std_logic_vector(7 downto 0);
    signal expr_193_wire_constant : std_logic_vector(2 downto 0);
    signal next_I_186 : std_logic_vector(2 downto 0);
    signal simple_obj_ref_187_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_187_scaled : std_logic_vector(2 downto 0);
    signal type_cast_179_wire_constant : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    array_obj_ref_188_offset_scale_factor_0 <= "001";
    array_obj_ref_188_resized_base_address <= "000";
    array_obj_ref_188_word_offset_0 <= "000";
    expr_184_wire_constant <= "001";
    expr_189_wire_constant <= "00000000";
    expr_193_wire_constant <= "100";
    type_cast_179_wire_constant <= "000";
    phi_stmt_175: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_179_wire_constant & next_I_186;
      req <= phi_stmt_175_req_0 & phi_stmt_175_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_175_ack_0,
          idata => idata,
          odata => I_0_175,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_175
    array_obj_ref_188_index_0_resize: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => I_0_175, dout => simple_obj_ref_187_resized, req => array_obj_ref_188_index_0_resize_req_0, ack => array_obj_ref_188_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_188_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_187_scaled, dout => array_obj_ref_188_final_offset, req => array_obj_ref_188_offset_inst_req_0, ack => array_obj_ref_188_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_188_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_188_addr_0_ack_0 <= array_obj_ref_188_addr_0_req_0;
      aggregated_sig <= array_obj_ref_188_root_address;
      array_obj_ref_188_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_188_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_188_gather_scatter_ack_0 <= array_obj_ref_188_gather_scatter_req_0;
      aggregated_sig <= expr_189_wire_constant;
      array_obj_ref_188_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_188_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_188_index_0_rename_ack_0 <= array_obj_ref_188_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_187_resized;
      simple_obj_ref_187_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_188_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_188_root_address_inst_ack_0 <= array_obj_ref_188_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_188_final_offset;
      array_obj_ref_188_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    if_stmt_191_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_194_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_191_branch_req_0,
          ack0 => if_stmt_191_branch_ack_0,
          ack1 => if_stmt_191_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_185_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_0_175;
      next_I_186 <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "001",
          constant_width => 3,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_185_inst_req_0,
          ackL => binary_185_inst_ack_0,
          reqR => binary_185_inst_req_1,
          ackR => binary_185_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_194_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= next_I_186;
      binary_194_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "100",
          constant_width => 3,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_194_inst_req_0,
          ackL => binary_194_inst_ack_0,
          reqR => binary_194_inst_req_1,
          ackR => binary_194_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_188_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_188_store_0_req_0;
      array_obj_ref_188_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_188_store_0_req_1;
      array_obj_ref_188_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_188_word_address_0;
      data_in <= array_obj_ref_188_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(2 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_free_queue_ram is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_free_queue_ram;
architecture Default of default_initializer_free_queue_ram is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_free_queue_ram_CP_485_start: Boolean;
  -- links between control-path and data-path
  signal binary_214_inst_req_0 : boolean;
  signal binary_214_inst_ack_0 : boolean;
  signal binary_214_inst_req_1 : boolean;
  signal binary_214_inst_ack_1 : boolean;
  signal array_obj_ref_217_index_0_resize_req_0 : boolean;
  signal array_obj_ref_217_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_217_index_0_rename_req_0 : boolean;
  signal array_obj_ref_217_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_217_offset_inst_req_0 : boolean;
  signal array_obj_ref_217_offset_inst_ack_0 : boolean;
  signal array_obj_ref_217_root_address_inst_req_0 : boolean;
  signal array_obj_ref_217_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_217_root_address_inst_req_1 : boolean;
  signal array_obj_ref_217_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_217_addr_0_req_0 : boolean;
  signal array_obj_ref_217_addr_0_ack_0 : boolean;
  signal array_obj_ref_217_gather_scatter_req_0 : boolean;
  signal array_obj_ref_217_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_217_store_0_req_0 : boolean;
  signal array_obj_ref_217_store_0_ack_0 : boolean;
  signal array_obj_ref_217_store_0_req_1 : boolean;
  signal array_obj_ref_217_store_0_ack_1 : boolean;
  signal binary_223_inst_req_0 : boolean;
  signal binary_223_inst_ack_0 : boolean;
  signal binary_223_inst_req_1 : boolean;
  signal binary_223_inst_ack_1 : boolean;
  signal if_stmt_220_branch_req_0 : boolean;
  signal if_stmt_220_branch_ack_1 : boolean;
  signal if_stmt_220_branch_ack_0 : boolean;
  signal phi_stmt_204_req_0 : boolean;
  signal phi_stmt_204_req_1 : boolean;
  signal phi_stmt_204_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_free_queue_ram_CP_485: Block -- control-path 
    signal cp_elements: BooleanArray(31 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(27) & cp_elements(31));
    binary_214_inst_req_0 <= cp_elements(1);
    cp_elements(2) <= OrReduce(cp_elements(16) & cp_elements(24));
    cp_elements(3) <= binary_214_inst_ack_0;
    binary_214_inst_req_1 <= cp_elements(3);
    cp_elements(4) <= binary_214_inst_ack_1;
    array_obj_ref_217_index_0_resize_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_217_index_0_resize_ack_0;
    array_obj_ref_217_index_0_rename_req_0 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_217_index_0_rename_ack_0;
    array_obj_ref_217_offset_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_217_offset_inst_ack_0;
    array_obj_ref_217_root_address_inst_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_217_root_address_inst_ack_0;
    array_obj_ref_217_root_address_inst_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_217_root_address_inst_ack_1;
    array_obj_ref_217_addr_0_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_217_addr_0_ack_0;
    array_obj_ref_217_gather_scatter_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_217_gather_scatter_ack_0;
    array_obj_ref_217_store_0_req_0 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_217_store_0_ack_0;
    array_obj_ref_217_store_0_req_1 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_217_store_0_ack_1;
    cp_elements(14) <= cp_elements(13);
    cp_elements(15) <= false;
    cp_elements(16) <= cp_elements(15);
    cp_elements(17) <= cp_elements(13);
    binary_223_inst_req_0 <= cp_elements(17);
    cp_elements(18) <= binary_223_inst_ack_0;
    binary_223_inst_req_1 <= cp_elements(18);
    cp_elements(19) <= binary_223_inst_ack_1;
    if_stmt_220_branch_req_0 <= cp_elements(19);
    cp_elements(20) <= cp_elements(19);
    cp_elements(21) <= cp_elements(20);
    cp_elements(22) <= if_stmt_220_branch_ack_1;
    phi_stmt_204_req_1 <= cp_elements(22);
    cp_elements(23) <= cp_elements(20);
    cp_elements(24) <= if_stmt_220_branch_ack_0;
    cp_elements(25) <= cp_elements(0);
    cp_elements(26) <= false;
    cp_elements(27) <= cp_elements(26);
    cp_elements(28) <= cp_elements(0);
    phi_stmt_204_req_0 <= cp_elements(28);
    cp_elements(29) <= OrReduce(cp_elements(22) & cp_elements(28));
    cp_elements(30) <= cp_elements(29);
    cp_elements(31) <= phi_stmt_204_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_0_204 : std_logic_vector(10 downto 0);
    signal array_obj_ref_217_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_217_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_217_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_217_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_217_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_217_word_address_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_217_word_offset_0 : std_logic_vector(10 downto 0);
    signal binary_223_wire : std_logic_vector(0 downto 0);
    signal expr_213_wire_constant : std_logic_vector(10 downto 0);
    signal expr_218_wire_constant : std_logic_vector(7 downto 0);
    signal expr_222_wire_constant : std_logic_vector(10 downto 0);
    signal next_I_215 : std_logic_vector(10 downto 0);
    signal simple_obj_ref_216_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_216_scaled : std_logic_vector(10 downto 0);
    signal type_cast_208_wire_constant : std_logic_vector(10 downto 0);
    -- 
  begin -- 
    array_obj_ref_217_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_217_resized_base_address <= "00000000001";
    array_obj_ref_217_word_offset_0 <= "00000000000";
    expr_213_wire_constant <= "00000000001";
    expr_218_wire_constant <= "00000000";
    expr_222_wire_constant <= "10000000000";
    type_cast_208_wire_constant <= "00000000000";
    phi_stmt_204: Block -- phi operator 
      signal idata: std_logic_vector(21 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_208_wire_constant & next_I_215;
      req <= phi_stmt_204_req_0 & phi_stmt_204_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 11) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_204_ack_0,
          idata => idata,
          odata => I_0_204,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_204
    array_obj_ref_217_index_0_resize: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => I_0_204, dout => simple_obj_ref_216_resized, req => array_obj_ref_217_index_0_resize_req_0, ack => array_obj_ref_217_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_217_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_216_scaled, dout => array_obj_ref_217_final_offset, req => array_obj_ref_217_offset_inst_req_0, ack => array_obj_ref_217_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_217_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_217_addr_0_ack_0 <= array_obj_ref_217_addr_0_req_0;
      aggregated_sig <= array_obj_ref_217_root_address;
      array_obj_ref_217_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_217_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_217_gather_scatter_ack_0 <= array_obj_ref_217_gather_scatter_req_0;
      aggregated_sig <= expr_218_wire_constant;
      array_obj_ref_217_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_217_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_217_index_0_rename_ack_0 <= array_obj_ref_217_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_216_resized;
      simple_obj_ref_216_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    if_stmt_220_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_223_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_220_branch_req_0,
          ack0 => if_stmt_220_branch_ack_0,
          ack1 => if_stmt_220_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_217_root_address_inst binary_214_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_217_final_offset & I_0_204;
      array_obj_ref_217_root_address <= data_out(21 downto 11);
      next_I_215 <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_217_root_address_inst_req_0;
      reqL(0) <= binary_214_inst_req_0;
      array_obj_ref_217_root_address_inst_ack_0 <= ackL(1);
      binary_214_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_217_root_address_inst_req_1;
      reqR(0) <= binary_214_inst_req_1;
      array_obj_ref_217_root_address_inst_ack_1 <= ackR(1);
      binary_214_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_223_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= next_I_215;
      binary_223_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10000000000",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_223_inst_req_0,
          ackL => binary_223_inst_ack_0,
          reqR => binary_223_inst_req_1,
          ackR => binary_223_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_217_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_217_store_0_req_0;
      array_obj_ref_217_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_217_store_0_req_1;
      array_obj_ref_217_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_217_word_address_0;
      data_in <= array_obj_ref_217_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(10 downto 0),
          mdata => memory_space_0_sr_data(7 downto 0),
          mtag => memory_space_0_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(4 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr;
architecture Default of default_initializer_xx_xstr is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr_CP_621_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_284_gather_scatter_req_0 : boolean;
  signal array_obj_ref_264_store_0_ack_0 : boolean;
  signal array_obj_ref_264_store_0_req_0 : boolean;
  signal array_obj_ref_244_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_288_store_0_req_1 : boolean;
  signal array_obj_ref_240_store_0_req_0 : boolean;
  signal array_obj_ref_288_store_0_req_0 : boolean;
  signal array_obj_ref_244_store_0_req_0 : boolean;
  signal array_obj_ref_280_store_0_ack_1 : boolean;
  signal array_obj_ref_256_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_256_gather_scatter_req_0 : boolean;
  signal array_obj_ref_280_store_0_req_1 : boolean;
  signal array_obj_ref_240_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_296_store_0_req_0 : boolean;
  signal array_obj_ref_280_store_0_ack_0 : boolean;
  signal array_obj_ref_240_gather_scatter_req_0 : boolean;
  signal array_obj_ref_304_store_0_ack_0 : boolean;
  signal array_obj_ref_280_store_0_req_0 : boolean;
  signal array_obj_ref_304_store_0_req_0 : boolean;
  signal array_obj_ref_264_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_256_store_0_ack_1 : boolean;
  signal array_obj_ref_244_gather_scatter_req_0 : boolean;
  signal array_obj_ref_252_store_0_ack_1 : boolean;
  signal array_obj_ref_252_store_0_req_1 : boolean;
  signal array_obj_ref_252_store_0_ack_0 : boolean;
  signal array_obj_ref_252_store_0_req_0 : boolean;
  signal array_obj_ref_264_gather_scatter_req_0 : boolean;
  signal array_obj_ref_280_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_280_gather_scatter_req_0 : boolean;
  signal array_obj_ref_236_store_0_ack_1 : boolean;
  signal array_obj_ref_236_store_0_req_1 : boolean;
  signal array_obj_ref_236_store_0_ack_0 : boolean;
  signal array_obj_ref_296_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_236_store_0_req_0 : boolean;
  signal array_obj_ref_292_store_0_req_0 : boolean;
  signal array_obj_ref_284_store_0_ack_1 : boolean;
  signal array_obj_ref_300_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_296_gather_scatter_req_0 : boolean;
  signal array_obj_ref_284_store_0_req_1 : boolean;
  signal array_obj_ref_236_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_292_store_0_ack_0 : boolean;
  signal array_obj_ref_288_store_0_ack_0 : boolean;
  signal array_obj_ref_236_gather_scatter_req_0 : boolean;
  signal array_obj_ref_276_store_0_ack_1 : boolean;
  signal array_obj_ref_256_store_0_req_1 : boolean;
  signal array_obj_ref_288_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_304_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_300_gather_scatter_req_0 : boolean;
  signal array_obj_ref_244_store_0_req_1 : boolean;
  signal array_obj_ref_240_store_0_ack_1 : boolean;
  signal array_obj_ref_244_store_0_ack_0 : boolean;
  signal array_obj_ref_276_store_0_req_1 : boolean;
  signal array_obj_ref_276_store_0_ack_0 : boolean;
  signal array_obj_ref_296_store_0_ack_1 : boolean;
  signal array_obj_ref_260_store_0_ack_1 : boolean;
  signal array_obj_ref_252_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_276_store_0_req_0 : boolean;
  signal array_obj_ref_276_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_232_store_0_ack_1 : boolean;
  signal array_obj_ref_276_gather_scatter_req_0 : boolean;
  signal array_obj_ref_232_store_0_req_1 : boolean;
  signal array_obj_ref_284_store_0_ack_0 : boolean;
  signal array_obj_ref_260_store_0_req_1 : boolean;
  signal array_obj_ref_232_store_0_ack_0 : boolean;
  signal array_obj_ref_232_store_0_req_0 : boolean;
  signal array_obj_ref_260_store_0_ack_0 : boolean;
  signal array_obj_ref_252_gather_scatter_req_0 : boolean;
  signal array_obj_ref_284_store_0_req_0 : boolean;
  signal array_obj_ref_304_gather_scatter_req_0 : boolean;
  signal array_obj_ref_292_gather_scatter_req_0 : boolean;
  signal array_obj_ref_264_store_0_ack_1 : boolean;
  signal array_obj_ref_272_store_0_ack_1 : boolean;
  signal array_obj_ref_300_store_0_ack_1 : boolean;
  signal array_obj_ref_240_store_0_req_1 : boolean;
  signal array_obj_ref_232_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_272_store_0_req_1 : boolean;
  signal array_obj_ref_296_store_0_req_1 : boolean;
  signal array_obj_ref_260_store_0_req_0 : boolean;
  signal array_obj_ref_256_store_0_ack_0 : boolean;
  signal array_obj_ref_292_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_272_store_0_ack_0 : boolean;
  signal array_obj_ref_232_gather_scatter_req_0 : boolean;
  signal array_obj_ref_272_store_0_req_0 : boolean;
  signal array_obj_ref_272_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_272_gather_scatter_req_0 : boolean;
  signal array_obj_ref_292_store_0_ack_1 : boolean;
  signal array_obj_ref_248_store_0_ack_1 : boolean;
  signal array_obj_ref_248_store_0_req_1 : boolean;
  signal array_obj_ref_300_store_0_req_1 : boolean;
  signal array_obj_ref_288_gather_scatter_req_0 : boolean;
  signal array_obj_ref_300_store_0_ack_0 : boolean;
  signal array_obj_ref_304_store_0_ack_1 : boolean;
  signal array_obj_ref_248_store_0_ack_0 : boolean;
  signal array_obj_ref_248_store_0_req_0 : boolean;
  signal array_obj_ref_240_store_0_ack_0 : boolean;
  signal array_obj_ref_268_store_0_ack_1 : boolean;
  signal array_obj_ref_296_store_0_ack_0 : boolean;
  signal array_obj_ref_256_store_0_req_0 : boolean;
  signal array_obj_ref_268_store_0_req_1 : boolean;
  signal array_obj_ref_268_store_0_ack_0 : boolean;
  signal array_obj_ref_268_store_0_req_0 : boolean;
  signal array_obj_ref_268_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_288_store_0_ack_1 : boolean;
  signal array_obj_ref_260_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_268_gather_scatter_req_0 : boolean;
  signal array_obj_ref_292_store_0_req_1 : boolean;
  signal array_obj_ref_260_gather_scatter_req_0 : boolean;
  signal array_obj_ref_248_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_284_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_264_store_0_req_1 : boolean;
  signal array_obj_ref_248_gather_scatter_req_0 : boolean;
  signal array_obj_ref_300_store_0_req_0 : boolean;
  signal array_obj_ref_304_store_0_req_1 : boolean;
  signal array_obj_ref_244_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 19 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr_CP_621: Block -- control-path 
    signal cp_elements: BooleanArray(57 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(57);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(57), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_232_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_232_gather_scatter_ack_0;
    array_obj_ref_232_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_232_store_0_ack_0;
    array_obj_ref_232_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_232_store_0_ack_1;
    array_obj_ref_236_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_236_gather_scatter_ack_0;
    array_obj_ref_236_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_236_store_0_ack_0;
    array_obj_ref_236_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_236_store_0_ack_1;
    array_obj_ref_240_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_240_gather_scatter_ack_0;
    array_obj_ref_240_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_240_store_0_ack_0;
    array_obj_ref_240_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_240_store_0_ack_1;
    array_obj_ref_244_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_244_gather_scatter_ack_0;
    array_obj_ref_244_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_244_store_0_ack_0;
    array_obj_ref_244_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_244_store_0_ack_1;
    array_obj_ref_248_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_248_gather_scatter_ack_0;
    array_obj_ref_248_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_248_store_0_ack_0;
    array_obj_ref_248_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_248_store_0_ack_1;
    array_obj_ref_252_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_252_gather_scatter_ack_0;
    array_obj_ref_252_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_252_store_0_ack_0;
    array_obj_ref_252_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_252_store_0_ack_1;
    array_obj_ref_256_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_256_gather_scatter_ack_0;
    array_obj_ref_256_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_256_store_0_ack_0;
    array_obj_ref_256_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_256_store_0_ack_1;
    array_obj_ref_260_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_260_gather_scatter_ack_0;
    array_obj_ref_260_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_260_store_0_ack_0;
    array_obj_ref_260_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_260_store_0_ack_1;
    array_obj_ref_264_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_264_gather_scatter_ack_0;
    array_obj_ref_264_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_264_store_0_ack_0;
    array_obj_ref_264_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_264_store_0_ack_1;
    array_obj_ref_268_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_268_gather_scatter_ack_0;
    array_obj_ref_268_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_268_store_0_ack_0;
    array_obj_ref_268_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_268_store_0_ack_1;
    array_obj_ref_272_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_272_gather_scatter_ack_0;
    array_obj_ref_272_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_272_store_0_ack_0;
    array_obj_ref_272_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_272_store_0_ack_1;
    array_obj_ref_276_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_276_gather_scatter_ack_0;
    array_obj_ref_276_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_276_store_0_ack_0;
    array_obj_ref_276_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_276_store_0_ack_1;
    array_obj_ref_280_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_280_gather_scatter_ack_0;
    array_obj_ref_280_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_280_store_0_ack_0;
    array_obj_ref_280_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_280_store_0_ack_1;
    array_obj_ref_284_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_284_gather_scatter_ack_0;
    array_obj_ref_284_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_284_store_0_ack_0;
    array_obj_ref_284_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_284_store_0_ack_1;
    array_obj_ref_288_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_288_gather_scatter_ack_0;
    array_obj_ref_288_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_288_store_0_ack_0;
    array_obj_ref_288_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_288_store_0_ack_1;
    array_obj_ref_292_gather_scatter_req_0 <= cp_elements(45);
    cp_elements(46) <= array_obj_ref_292_gather_scatter_ack_0;
    array_obj_ref_292_store_0_req_0 <= cp_elements(46);
    cp_elements(47) <= array_obj_ref_292_store_0_ack_0;
    array_obj_ref_292_store_0_req_1 <= cp_elements(47);
    cp_elements(48) <= array_obj_ref_292_store_0_ack_1;
    array_obj_ref_296_gather_scatter_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_296_gather_scatter_ack_0;
    array_obj_ref_296_store_0_req_0 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_296_store_0_ack_0;
    array_obj_ref_296_store_0_req_1 <= cp_elements(50);
    cp_elements(51) <= array_obj_ref_296_store_0_ack_1;
    array_obj_ref_300_gather_scatter_req_0 <= cp_elements(51);
    cp_elements(52) <= array_obj_ref_300_gather_scatter_ack_0;
    array_obj_ref_300_store_0_req_0 <= cp_elements(52);
    cp_elements(53) <= array_obj_ref_300_store_0_ack_0;
    array_obj_ref_300_store_0_req_1 <= cp_elements(53);
    cp_elements(54) <= array_obj_ref_300_store_0_ack_1;
    array_obj_ref_304_gather_scatter_req_0 <= cp_elements(54);
    cp_elements(55) <= array_obj_ref_304_gather_scatter_ack_0;
    array_obj_ref_304_store_0_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_304_store_0_ack_0;
    array_obj_ref_304_store_0_req_1 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_304_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_232_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_232_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_236_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_236_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_240_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_240_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_244_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_244_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_248_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_248_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_252_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_252_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_256_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_256_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_260_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_260_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_264_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_264_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_268_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_268_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_272_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_272_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_276_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_276_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_280_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_280_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_284_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_284_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_288_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_288_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_292_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_292_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_296_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_296_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_300_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_300_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_304_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_304_word_address_0 : std_logic_vector(4 downto 0);
    signal expr_233_wire_constant : std_logic_vector(7 downto 0);
    signal expr_237_wire_constant : std_logic_vector(7 downto 0);
    signal expr_241_wire_constant : std_logic_vector(7 downto 0);
    signal expr_245_wire_constant : std_logic_vector(7 downto 0);
    signal expr_249_wire_constant : std_logic_vector(7 downto 0);
    signal expr_253_wire_constant : std_logic_vector(7 downto 0);
    signal expr_257_wire_constant : std_logic_vector(7 downto 0);
    signal expr_261_wire_constant : std_logic_vector(7 downto 0);
    signal expr_265_wire_constant : std_logic_vector(7 downto 0);
    signal expr_269_wire_constant : std_logic_vector(7 downto 0);
    signal expr_273_wire_constant : std_logic_vector(7 downto 0);
    signal expr_277_wire_constant : std_logic_vector(7 downto 0);
    signal expr_281_wire_constant : std_logic_vector(7 downto 0);
    signal expr_285_wire_constant : std_logic_vector(7 downto 0);
    signal expr_289_wire_constant : std_logic_vector(7 downto 0);
    signal expr_293_wire_constant : std_logic_vector(7 downto 0);
    signal expr_297_wire_constant : std_logic_vector(7 downto 0);
    signal expr_301_wire_constant : std_logic_vector(7 downto 0);
    signal expr_305_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_232_word_address_0 <= "00000";
    array_obj_ref_236_word_address_0 <= "00001";
    array_obj_ref_240_word_address_0 <= "00010";
    array_obj_ref_244_word_address_0 <= "00011";
    array_obj_ref_248_word_address_0 <= "00100";
    array_obj_ref_252_word_address_0 <= "00101";
    array_obj_ref_256_word_address_0 <= "00110";
    array_obj_ref_260_word_address_0 <= "00111";
    array_obj_ref_264_word_address_0 <= "01000";
    array_obj_ref_268_word_address_0 <= "01001";
    array_obj_ref_272_word_address_0 <= "01010";
    array_obj_ref_276_word_address_0 <= "01011";
    array_obj_ref_280_word_address_0 <= "01100";
    array_obj_ref_284_word_address_0 <= "01101";
    array_obj_ref_288_word_address_0 <= "01110";
    array_obj_ref_292_word_address_0 <= "01111";
    array_obj_ref_296_word_address_0 <= "10000";
    array_obj_ref_300_word_address_0 <= "10001";
    array_obj_ref_304_word_address_0 <= "10010";
    expr_233_wire_constant <= "01100110";
    expr_237_wire_constant <= "01110010";
    expr_241_wire_constant <= "01100101";
    expr_245_wire_constant <= "01100101";
    expr_249_wire_constant <= "01011111";
    expr_253_wire_constant <= "01110001";
    expr_257_wire_constant <= "01110101";
    expr_261_wire_constant <= "01100101";
    expr_265_wire_constant <= "01110101";
    expr_269_wire_constant <= "01100101";
    expr_273_wire_constant <= "01011111";
    expr_277_wire_constant <= "01110010";
    expr_281_wire_constant <= "01100101";
    expr_285_wire_constant <= "01110001";
    expr_289_wire_constant <= "01110101";
    expr_293_wire_constant <= "01100101";
    expr_297_wire_constant <= "01110011";
    expr_301_wire_constant <= "01110100";
    expr_305_wire_constant <= "00000000";
    array_obj_ref_232_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_232_gather_scatter_ack_0 <= array_obj_ref_232_gather_scatter_req_0;
      aggregated_sig <= expr_233_wire_constant;
      array_obj_ref_232_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_236_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_236_gather_scatter_ack_0 <= array_obj_ref_236_gather_scatter_req_0;
      aggregated_sig <= expr_237_wire_constant;
      array_obj_ref_236_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_240_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_240_gather_scatter_ack_0 <= array_obj_ref_240_gather_scatter_req_0;
      aggregated_sig <= expr_241_wire_constant;
      array_obj_ref_240_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_244_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_244_gather_scatter_ack_0 <= array_obj_ref_244_gather_scatter_req_0;
      aggregated_sig <= expr_245_wire_constant;
      array_obj_ref_244_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_248_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_248_gather_scatter_ack_0 <= array_obj_ref_248_gather_scatter_req_0;
      aggregated_sig <= expr_249_wire_constant;
      array_obj_ref_248_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_252_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_252_gather_scatter_ack_0 <= array_obj_ref_252_gather_scatter_req_0;
      aggregated_sig <= expr_253_wire_constant;
      array_obj_ref_252_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_256_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_256_gather_scatter_ack_0 <= array_obj_ref_256_gather_scatter_req_0;
      aggregated_sig <= expr_257_wire_constant;
      array_obj_ref_256_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_260_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_260_gather_scatter_ack_0 <= array_obj_ref_260_gather_scatter_req_0;
      aggregated_sig <= expr_261_wire_constant;
      array_obj_ref_260_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_264_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_264_gather_scatter_ack_0 <= array_obj_ref_264_gather_scatter_req_0;
      aggregated_sig <= expr_265_wire_constant;
      array_obj_ref_264_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_268_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_268_gather_scatter_ack_0 <= array_obj_ref_268_gather_scatter_req_0;
      aggregated_sig <= expr_269_wire_constant;
      array_obj_ref_268_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_272_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_272_gather_scatter_ack_0 <= array_obj_ref_272_gather_scatter_req_0;
      aggregated_sig <= expr_273_wire_constant;
      array_obj_ref_272_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_276_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_276_gather_scatter_ack_0 <= array_obj_ref_276_gather_scatter_req_0;
      aggregated_sig <= expr_277_wire_constant;
      array_obj_ref_276_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_280_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_280_gather_scatter_ack_0 <= array_obj_ref_280_gather_scatter_req_0;
      aggregated_sig <= expr_281_wire_constant;
      array_obj_ref_280_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_284_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_284_gather_scatter_ack_0 <= array_obj_ref_284_gather_scatter_req_0;
      aggregated_sig <= expr_285_wire_constant;
      array_obj_ref_284_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_288_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_288_gather_scatter_ack_0 <= array_obj_ref_288_gather_scatter_req_0;
      aggregated_sig <= expr_289_wire_constant;
      array_obj_ref_288_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_292_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_292_gather_scatter_ack_0 <= array_obj_ref_292_gather_scatter_req_0;
      aggregated_sig <= expr_293_wire_constant;
      array_obj_ref_292_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_296_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_296_gather_scatter_ack_0 <= array_obj_ref_296_gather_scatter_req_0;
      aggregated_sig <= expr_297_wire_constant;
      array_obj_ref_296_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_300_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_300_gather_scatter_ack_0 <= array_obj_ref_300_gather_scatter_req_0;
      aggregated_sig <= expr_301_wire_constant;
      array_obj_ref_300_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_304_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_304_gather_scatter_ack_0 <= array_obj_ref_304_gather_scatter_req_0;
      aggregated_sig <= expr_305_wire_constant;
      array_obj_ref_304_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_244_store_0 array_obj_ref_240_store_0 array_obj_ref_256_store_0 array_obj_ref_232_store_0 array_obj_ref_236_store_0 array_obj_ref_268_store_0 array_obj_ref_288_store_0 array_obj_ref_284_store_0 array_obj_ref_300_store_0 array_obj_ref_292_store_0 array_obj_ref_280_store_0 array_obj_ref_276_store_0 array_obj_ref_252_store_0 array_obj_ref_248_store_0 array_obj_ref_304_store_0 array_obj_ref_264_store_0 array_obj_ref_260_store_0 array_obj_ref_272_store_0 array_obj_ref_296_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(94 downto 0);
      signal data_in: std_logic_vector(151 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 18 downto 0);
      -- 
    begin -- 
      reqL(18) <= array_obj_ref_244_store_0_req_0;
      reqL(17) <= array_obj_ref_240_store_0_req_0;
      reqL(16) <= array_obj_ref_256_store_0_req_0;
      reqL(15) <= array_obj_ref_232_store_0_req_0;
      reqL(14) <= array_obj_ref_236_store_0_req_0;
      reqL(13) <= array_obj_ref_268_store_0_req_0;
      reqL(12) <= array_obj_ref_288_store_0_req_0;
      reqL(11) <= array_obj_ref_284_store_0_req_0;
      reqL(10) <= array_obj_ref_300_store_0_req_0;
      reqL(9) <= array_obj_ref_292_store_0_req_0;
      reqL(8) <= array_obj_ref_280_store_0_req_0;
      reqL(7) <= array_obj_ref_276_store_0_req_0;
      reqL(6) <= array_obj_ref_252_store_0_req_0;
      reqL(5) <= array_obj_ref_248_store_0_req_0;
      reqL(4) <= array_obj_ref_304_store_0_req_0;
      reqL(3) <= array_obj_ref_264_store_0_req_0;
      reqL(2) <= array_obj_ref_260_store_0_req_0;
      reqL(1) <= array_obj_ref_272_store_0_req_0;
      reqL(0) <= array_obj_ref_296_store_0_req_0;
      array_obj_ref_244_store_0_ack_0 <= ackL(18);
      array_obj_ref_240_store_0_ack_0 <= ackL(17);
      array_obj_ref_256_store_0_ack_0 <= ackL(16);
      array_obj_ref_232_store_0_ack_0 <= ackL(15);
      array_obj_ref_236_store_0_ack_0 <= ackL(14);
      array_obj_ref_268_store_0_ack_0 <= ackL(13);
      array_obj_ref_288_store_0_ack_0 <= ackL(12);
      array_obj_ref_284_store_0_ack_0 <= ackL(11);
      array_obj_ref_300_store_0_ack_0 <= ackL(10);
      array_obj_ref_292_store_0_ack_0 <= ackL(9);
      array_obj_ref_280_store_0_ack_0 <= ackL(8);
      array_obj_ref_276_store_0_ack_0 <= ackL(7);
      array_obj_ref_252_store_0_ack_0 <= ackL(6);
      array_obj_ref_248_store_0_ack_0 <= ackL(5);
      array_obj_ref_304_store_0_ack_0 <= ackL(4);
      array_obj_ref_264_store_0_ack_0 <= ackL(3);
      array_obj_ref_260_store_0_ack_0 <= ackL(2);
      array_obj_ref_272_store_0_ack_0 <= ackL(1);
      array_obj_ref_296_store_0_ack_0 <= ackL(0);
      reqR(18) <= array_obj_ref_244_store_0_req_1;
      reqR(17) <= array_obj_ref_240_store_0_req_1;
      reqR(16) <= array_obj_ref_256_store_0_req_1;
      reqR(15) <= array_obj_ref_232_store_0_req_1;
      reqR(14) <= array_obj_ref_236_store_0_req_1;
      reqR(13) <= array_obj_ref_268_store_0_req_1;
      reqR(12) <= array_obj_ref_288_store_0_req_1;
      reqR(11) <= array_obj_ref_284_store_0_req_1;
      reqR(10) <= array_obj_ref_300_store_0_req_1;
      reqR(9) <= array_obj_ref_292_store_0_req_1;
      reqR(8) <= array_obj_ref_280_store_0_req_1;
      reqR(7) <= array_obj_ref_276_store_0_req_1;
      reqR(6) <= array_obj_ref_252_store_0_req_1;
      reqR(5) <= array_obj_ref_248_store_0_req_1;
      reqR(4) <= array_obj_ref_304_store_0_req_1;
      reqR(3) <= array_obj_ref_264_store_0_req_1;
      reqR(2) <= array_obj_ref_260_store_0_req_1;
      reqR(1) <= array_obj_ref_272_store_0_req_1;
      reqR(0) <= array_obj_ref_296_store_0_req_1;
      array_obj_ref_244_store_0_ack_1 <= ackR(18);
      array_obj_ref_240_store_0_ack_1 <= ackR(17);
      array_obj_ref_256_store_0_ack_1 <= ackR(16);
      array_obj_ref_232_store_0_ack_1 <= ackR(15);
      array_obj_ref_236_store_0_ack_1 <= ackR(14);
      array_obj_ref_268_store_0_ack_1 <= ackR(13);
      array_obj_ref_288_store_0_ack_1 <= ackR(12);
      array_obj_ref_284_store_0_ack_1 <= ackR(11);
      array_obj_ref_300_store_0_ack_1 <= ackR(10);
      array_obj_ref_292_store_0_ack_1 <= ackR(9);
      array_obj_ref_280_store_0_ack_1 <= ackR(8);
      array_obj_ref_276_store_0_ack_1 <= ackR(7);
      array_obj_ref_252_store_0_ack_1 <= ackR(6);
      array_obj_ref_248_store_0_ack_1 <= ackR(5);
      array_obj_ref_304_store_0_ack_1 <= ackR(4);
      array_obj_ref_264_store_0_ack_1 <= ackR(3);
      array_obj_ref_260_store_0_ack_1 <= ackR(2);
      array_obj_ref_272_store_0_ack_1 <= ackR(1);
      array_obj_ref_296_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_244_word_address_0 & array_obj_ref_240_word_address_0 & array_obj_ref_256_word_address_0 & array_obj_ref_232_word_address_0 & array_obj_ref_236_word_address_0 & array_obj_ref_268_word_address_0 & array_obj_ref_288_word_address_0 & array_obj_ref_284_word_address_0 & array_obj_ref_300_word_address_0 & array_obj_ref_292_word_address_0 & array_obj_ref_280_word_address_0 & array_obj_ref_276_word_address_0 & array_obj_ref_252_word_address_0 & array_obj_ref_248_word_address_0 & array_obj_ref_304_word_address_0 & array_obj_ref_264_word_address_0 & array_obj_ref_260_word_address_0 & array_obj_ref_272_word_address_0 & array_obj_ref_296_word_address_0;
      data_in <= array_obj_ref_244_data_0 & array_obj_ref_240_data_0 & array_obj_ref_256_data_0 & array_obj_ref_232_data_0 & array_obj_ref_236_data_0 & array_obj_ref_268_data_0 & array_obj_ref_288_data_0 & array_obj_ref_284_data_0 & array_obj_ref_300_data_0 & array_obj_ref_292_data_0 & array_obj_ref_280_data_0 & array_obj_ref_276_data_0 & array_obj_ref_252_data_0 & array_obj_ref_248_data_0 & array_obj_ref_304_data_0 & array_obj_ref_264_data_0 & array_obj_ref_260_data_0 & array_obj_ref_272_data_0 & array_obj_ref_296_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 5,
        data_width => 8,
        num_reqs => 19,
        tag_length => 5,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(4 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 19,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr1;
architecture Default of default_initializer_xx_xstr1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr1_CP_1023_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_310_gather_scatter_req_0 : boolean;
  signal array_obj_ref_310_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_310_store_0_req_0 : boolean;
  signal array_obj_ref_310_store_0_ack_0 : boolean;
  signal array_obj_ref_310_store_0_req_1 : boolean;
  signal array_obj_ref_310_store_0_ack_1 : boolean;
  signal array_obj_ref_314_gather_scatter_req_0 : boolean;
  signal array_obj_ref_314_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_314_store_0_req_0 : boolean;
  signal array_obj_ref_314_store_0_ack_0 : boolean;
  signal array_obj_ref_314_store_0_req_1 : boolean;
  signal array_obj_ref_314_store_0_ack_1 : boolean;
  signal array_obj_ref_318_gather_scatter_req_0 : boolean;
  signal array_obj_ref_318_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_0 : boolean;
  signal array_obj_ref_318_store_0_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_1 : boolean;
  signal array_obj_ref_318_store_0_ack_1 : boolean;
  signal array_obj_ref_322_gather_scatter_req_0 : boolean;
  signal array_obj_ref_322_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_322_store_0_req_0 : boolean;
  signal array_obj_ref_322_store_0_ack_0 : boolean;
  signal array_obj_ref_322_store_0_req_1 : boolean;
  signal array_obj_ref_322_store_0_ack_1 : boolean;
  signal array_obj_ref_326_gather_scatter_req_0 : boolean;
  signal array_obj_ref_326_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_326_store_0_req_0 : boolean;
  signal array_obj_ref_326_store_0_ack_0 : boolean;
  signal array_obj_ref_326_store_0_req_1 : boolean;
  signal array_obj_ref_326_store_0_ack_1 : boolean;
  signal array_obj_ref_330_gather_scatter_req_0 : boolean;
  signal array_obj_ref_330_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_330_store_0_req_0 : boolean;
  signal array_obj_ref_330_store_0_ack_0 : boolean;
  signal array_obj_ref_330_store_0_req_1 : boolean;
  signal array_obj_ref_330_store_0_ack_1 : boolean;
  signal array_obj_ref_334_gather_scatter_req_0 : boolean;
  signal array_obj_ref_334_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_334_store_0_req_0 : boolean;
  signal array_obj_ref_334_store_0_ack_0 : boolean;
  signal array_obj_ref_334_store_0_req_1 : boolean;
  signal array_obj_ref_334_store_0_ack_1 : boolean;
  signal array_obj_ref_338_gather_scatter_req_0 : boolean;
  signal array_obj_ref_338_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_338_store_0_req_0 : boolean;
  signal array_obj_ref_338_store_0_ack_0 : boolean;
  signal array_obj_ref_338_store_0_req_1 : boolean;
  signal array_obj_ref_338_store_0_ack_1 : boolean;
  signal array_obj_ref_342_gather_scatter_req_0 : boolean;
  signal array_obj_ref_342_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_342_store_0_req_0 : boolean;
  signal array_obj_ref_342_store_0_ack_0 : boolean;
  signal array_obj_ref_342_store_0_req_1 : boolean;
  signal array_obj_ref_342_store_0_ack_1 : boolean;
  signal array_obj_ref_346_gather_scatter_req_0 : boolean;
  signal array_obj_ref_346_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_0 : boolean;
  signal array_obj_ref_346_store_0_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_1 : boolean;
  signal array_obj_ref_346_store_0_ack_1 : boolean;
  signal array_obj_ref_350_gather_scatter_req_0 : boolean;
  signal array_obj_ref_350_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_350_store_0_req_0 : boolean;
  signal array_obj_ref_350_store_0_ack_0 : boolean;
  signal array_obj_ref_350_store_0_req_1 : boolean;
  signal array_obj_ref_350_store_0_ack_1 : boolean;
  signal array_obj_ref_354_gather_scatter_req_0 : boolean;
  signal array_obj_ref_354_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_354_store_0_req_0 : boolean;
  signal array_obj_ref_354_store_0_ack_0 : boolean;
  signal array_obj_ref_354_store_0_req_1 : boolean;
  signal array_obj_ref_354_store_0_ack_1 : boolean;
  signal array_obj_ref_358_gather_scatter_req_0 : boolean;
  signal array_obj_ref_358_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_358_store_0_req_0 : boolean;
  signal array_obj_ref_358_store_0_ack_0 : boolean;
  signal array_obj_ref_358_store_0_req_1 : boolean;
  signal array_obj_ref_358_store_0_ack_1 : boolean;
  signal array_obj_ref_362_gather_scatter_req_0 : boolean;
  signal array_obj_ref_362_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_362_store_0_req_0 : boolean;
  signal array_obj_ref_362_store_0_ack_0 : boolean;
  signal array_obj_ref_362_store_0_req_1 : boolean;
  signal array_obj_ref_362_store_0_ack_1 : boolean;
  signal array_obj_ref_366_gather_scatter_req_0 : boolean;
  signal array_obj_ref_366_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_366_store_0_req_0 : boolean;
  signal array_obj_ref_366_store_0_ack_0 : boolean;
  signal array_obj_ref_366_store_0_req_1 : boolean;
  signal array_obj_ref_366_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 15 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr1_CP_1023: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_310_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_310_gather_scatter_ack_0;
    array_obj_ref_310_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_310_store_0_ack_0;
    array_obj_ref_310_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_310_store_0_ack_1;
    array_obj_ref_314_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_314_gather_scatter_ack_0;
    array_obj_ref_314_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_314_store_0_ack_0;
    array_obj_ref_314_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_314_store_0_ack_1;
    array_obj_ref_318_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_318_gather_scatter_ack_0;
    array_obj_ref_318_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_318_store_0_ack_0;
    array_obj_ref_318_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_318_store_0_ack_1;
    array_obj_ref_322_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_322_gather_scatter_ack_0;
    array_obj_ref_322_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_322_store_0_ack_0;
    array_obj_ref_322_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_322_store_0_ack_1;
    array_obj_ref_326_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_326_gather_scatter_ack_0;
    array_obj_ref_326_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_326_store_0_ack_0;
    array_obj_ref_326_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_326_store_0_ack_1;
    array_obj_ref_330_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_330_gather_scatter_ack_0;
    array_obj_ref_330_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_330_store_0_ack_0;
    array_obj_ref_330_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_330_store_0_ack_1;
    array_obj_ref_334_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_334_gather_scatter_ack_0;
    array_obj_ref_334_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_334_store_0_ack_0;
    array_obj_ref_334_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_334_store_0_ack_1;
    array_obj_ref_338_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_338_gather_scatter_ack_0;
    array_obj_ref_338_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_338_store_0_ack_0;
    array_obj_ref_338_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_338_store_0_ack_1;
    array_obj_ref_342_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_342_gather_scatter_ack_0;
    array_obj_ref_342_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_342_store_0_ack_0;
    array_obj_ref_342_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_342_store_0_ack_1;
    array_obj_ref_346_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_346_gather_scatter_ack_0;
    array_obj_ref_346_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_346_store_0_ack_0;
    array_obj_ref_346_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_346_store_0_ack_1;
    array_obj_ref_350_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_350_gather_scatter_ack_0;
    array_obj_ref_350_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_350_store_0_ack_0;
    array_obj_ref_350_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_350_store_0_ack_1;
    array_obj_ref_354_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_354_gather_scatter_ack_0;
    array_obj_ref_354_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_354_store_0_ack_0;
    array_obj_ref_354_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_354_store_0_ack_1;
    array_obj_ref_358_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_358_gather_scatter_ack_0;
    array_obj_ref_358_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_358_store_0_ack_0;
    array_obj_ref_358_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_358_store_0_ack_1;
    array_obj_ref_362_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_362_gather_scatter_ack_0;
    array_obj_ref_362_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_362_store_0_ack_0;
    array_obj_ref_362_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_362_store_0_ack_1;
    array_obj_ref_366_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_366_gather_scatter_ack_0;
    array_obj_ref_366_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_366_store_0_ack_0;
    array_obj_ref_366_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_366_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_310_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_310_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_314_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_314_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_318_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_318_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_322_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_322_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_326_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_326_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_330_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_330_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_334_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_334_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_338_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_338_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_342_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_342_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_346_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_346_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_350_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_350_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_354_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_354_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_358_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_358_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_362_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_362_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_366_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_366_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_311_wire_constant : std_logic_vector(7 downto 0);
    signal expr_315_wire_constant : std_logic_vector(7 downto 0);
    signal expr_319_wire_constant : std_logic_vector(7 downto 0);
    signal expr_323_wire_constant : std_logic_vector(7 downto 0);
    signal expr_327_wire_constant : std_logic_vector(7 downto 0);
    signal expr_331_wire_constant : std_logic_vector(7 downto 0);
    signal expr_335_wire_constant : std_logic_vector(7 downto 0);
    signal expr_339_wire_constant : std_logic_vector(7 downto 0);
    signal expr_343_wire_constant : std_logic_vector(7 downto 0);
    signal expr_347_wire_constant : std_logic_vector(7 downto 0);
    signal expr_351_wire_constant : std_logic_vector(7 downto 0);
    signal expr_355_wire_constant : std_logic_vector(7 downto 0);
    signal expr_359_wire_constant : std_logic_vector(7 downto 0);
    signal expr_363_wire_constant : std_logic_vector(7 downto 0);
    signal expr_367_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_310_word_address_0 <= "0000";
    array_obj_ref_314_word_address_0 <= "0001";
    array_obj_ref_318_word_address_0 <= "0010";
    array_obj_ref_322_word_address_0 <= "0011";
    array_obj_ref_326_word_address_0 <= "0100";
    array_obj_ref_330_word_address_0 <= "0101";
    array_obj_ref_334_word_address_0 <= "0110";
    array_obj_ref_338_word_address_0 <= "0111";
    array_obj_ref_342_word_address_0 <= "1000";
    array_obj_ref_346_word_address_0 <= "1001";
    array_obj_ref_350_word_address_0 <= "1010";
    array_obj_ref_354_word_address_0 <= "1011";
    array_obj_ref_358_word_address_0 <= "1100";
    array_obj_ref_362_word_address_0 <= "1101";
    array_obj_ref_366_word_address_0 <= "1110";
    expr_311_wire_constant <= "01100110";
    expr_315_wire_constant <= "01110010";
    expr_319_wire_constant <= "01100101";
    expr_323_wire_constant <= "01100101";
    expr_327_wire_constant <= "01011111";
    expr_331_wire_constant <= "01110001";
    expr_335_wire_constant <= "01110101";
    expr_339_wire_constant <= "01100101";
    expr_343_wire_constant <= "01110101";
    expr_347_wire_constant <= "01100101";
    expr_351_wire_constant <= "01011111";
    expr_355_wire_constant <= "01100001";
    expr_359_wire_constant <= "01100011";
    expr_363_wire_constant <= "01101011";
    expr_367_wire_constant <= "00000000";
    array_obj_ref_310_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_310_gather_scatter_ack_0 <= array_obj_ref_310_gather_scatter_req_0;
      aggregated_sig <= expr_311_wire_constant;
      array_obj_ref_310_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_314_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_314_gather_scatter_ack_0 <= array_obj_ref_314_gather_scatter_req_0;
      aggregated_sig <= expr_315_wire_constant;
      array_obj_ref_314_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_318_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_318_gather_scatter_ack_0 <= array_obj_ref_318_gather_scatter_req_0;
      aggregated_sig <= expr_319_wire_constant;
      array_obj_ref_318_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_322_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_322_gather_scatter_ack_0 <= array_obj_ref_322_gather_scatter_req_0;
      aggregated_sig <= expr_323_wire_constant;
      array_obj_ref_322_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_326_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_326_gather_scatter_ack_0 <= array_obj_ref_326_gather_scatter_req_0;
      aggregated_sig <= expr_327_wire_constant;
      array_obj_ref_326_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_330_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_330_gather_scatter_ack_0 <= array_obj_ref_330_gather_scatter_req_0;
      aggregated_sig <= expr_331_wire_constant;
      array_obj_ref_330_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_334_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_334_gather_scatter_ack_0 <= array_obj_ref_334_gather_scatter_req_0;
      aggregated_sig <= expr_335_wire_constant;
      array_obj_ref_334_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_338_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_338_gather_scatter_ack_0 <= array_obj_ref_338_gather_scatter_req_0;
      aggregated_sig <= expr_339_wire_constant;
      array_obj_ref_338_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_342_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_342_gather_scatter_ack_0 <= array_obj_ref_342_gather_scatter_req_0;
      aggregated_sig <= expr_343_wire_constant;
      array_obj_ref_342_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_346_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_346_gather_scatter_ack_0 <= array_obj_ref_346_gather_scatter_req_0;
      aggregated_sig <= expr_347_wire_constant;
      array_obj_ref_346_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_350_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_350_gather_scatter_ack_0 <= array_obj_ref_350_gather_scatter_req_0;
      aggregated_sig <= expr_351_wire_constant;
      array_obj_ref_350_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_354_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_354_gather_scatter_ack_0 <= array_obj_ref_354_gather_scatter_req_0;
      aggregated_sig <= expr_355_wire_constant;
      array_obj_ref_354_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_358_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_358_gather_scatter_ack_0 <= array_obj_ref_358_gather_scatter_req_0;
      aggregated_sig <= expr_359_wire_constant;
      array_obj_ref_358_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_362_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_362_gather_scatter_ack_0 <= array_obj_ref_362_gather_scatter_req_0;
      aggregated_sig <= expr_363_wire_constant;
      array_obj_ref_362_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_366_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_366_gather_scatter_ack_0 <= array_obj_ref_366_gather_scatter_req_0;
      aggregated_sig <= expr_367_wire_constant;
      array_obj_ref_366_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_342_store_0 array_obj_ref_326_store_0 array_obj_ref_330_store_0 array_obj_ref_318_store_0 array_obj_ref_358_store_0 array_obj_ref_362_store_0 array_obj_ref_334_store_0 array_obj_ref_346_store_0 array_obj_ref_310_store_0 array_obj_ref_314_store_0 array_obj_ref_322_store_0 array_obj_ref_350_store_0 array_obj_ref_338_store_0 array_obj_ref_354_store_0 array_obj_ref_366_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(59 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_342_store_0_req_0;
      reqL(13) <= array_obj_ref_326_store_0_req_0;
      reqL(12) <= array_obj_ref_330_store_0_req_0;
      reqL(11) <= array_obj_ref_318_store_0_req_0;
      reqL(10) <= array_obj_ref_358_store_0_req_0;
      reqL(9) <= array_obj_ref_362_store_0_req_0;
      reqL(8) <= array_obj_ref_334_store_0_req_0;
      reqL(7) <= array_obj_ref_346_store_0_req_0;
      reqL(6) <= array_obj_ref_310_store_0_req_0;
      reqL(5) <= array_obj_ref_314_store_0_req_0;
      reqL(4) <= array_obj_ref_322_store_0_req_0;
      reqL(3) <= array_obj_ref_350_store_0_req_0;
      reqL(2) <= array_obj_ref_338_store_0_req_0;
      reqL(1) <= array_obj_ref_354_store_0_req_0;
      reqL(0) <= array_obj_ref_366_store_0_req_0;
      array_obj_ref_342_store_0_ack_0 <= ackL(14);
      array_obj_ref_326_store_0_ack_0 <= ackL(13);
      array_obj_ref_330_store_0_ack_0 <= ackL(12);
      array_obj_ref_318_store_0_ack_0 <= ackL(11);
      array_obj_ref_358_store_0_ack_0 <= ackL(10);
      array_obj_ref_362_store_0_ack_0 <= ackL(9);
      array_obj_ref_334_store_0_ack_0 <= ackL(8);
      array_obj_ref_346_store_0_ack_0 <= ackL(7);
      array_obj_ref_310_store_0_ack_0 <= ackL(6);
      array_obj_ref_314_store_0_ack_0 <= ackL(5);
      array_obj_ref_322_store_0_ack_0 <= ackL(4);
      array_obj_ref_350_store_0_ack_0 <= ackL(3);
      array_obj_ref_338_store_0_ack_0 <= ackL(2);
      array_obj_ref_354_store_0_ack_0 <= ackL(1);
      array_obj_ref_366_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_342_store_0_req_1;
      reqR(13) <= array_obj_ref_326_store_0_req_1;
      reqR(12) <= array_obj_ref_330_store_0_req_1;
      reqR(11) <= array_obj_ref_318_store_0_req_1;
      reqR(10) <= array_obj_ref_358_store_0_req_1;
      reqR(9) <= array_obj_ref_362_store_0_req_1;
      reqR(8) <= array_obj_ref_334_store_0_req_1;
      reqR(7) <= array_obj_ref_346_store_0_req_1;
      reqR(6) <= array_obj_ref_310_store_0_req_1;
      reqR(5) <= array_obj_ref_314_store_0_req_1;
      reqR(4) <= array_obj_ref_322_store_0_req_1;
      reqR(3) <= array_obj_ref_350_store_0_req_1;
      reqR(2) <= array_obj_ref_338_store_0_req_1;
      reqR(1) <= array_obj_ref_354_store_0_req_1;
      reqR(0) <= array_obj_ref_366_store_0_req_1;
      array_obj_ref_342_store_0_ack_1 <= ackR(14);
      array_obj_ref_326_store_0_ack_1 <= ackR(13);
      array_obj_ref_330_store_0_ack_1 <= ackR(12);
      array_obj_ref_318_store_0_ack_1 <= ackR(11);
      array_obj_ref_358_store_0_ack_1 <= ackR(10);
      array_obj_ref_362_store_0_ack_1 <= ackR(9);
      array_obj_ref_334_store_0_ack_1 <= ackR(8);
      array_obj_ref_346_store_0_ack_1 <= ackR(7);
      array_obj_ref_310_store_0_ack_1 <= ackR(6);
      array_obj_ref_314_store_0_ack_1 <= ackR(5);
      array_obj_ref_322_store_0_ack_1 <= ackR(4);
      array_obj_ref_350_store_0_ack_1 <= ackR(3);
      array_obj_ref_338_store_0_ack_1 <= ackR(2);
      array_obj_ref_354_store_0_ack_1 <= ackR(1);
      array_obj_ref_366_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_342_word_address_0 & array_obj_ref_326_word_address_0 & array_obj_ref_330_word_address_0 & array_obj_ref_318_word_address_0 & array_obj_ref_358_word_address_0 & array_obj_ref_362_word_address_0 & array_obj_ref_334_word_address_0 & array_obj_ref_346_word_address_0 & array_obj_ref_310_word_address_0 & array_obj_ref_314_word_address_0 & array_obj_ref_322_word_address_0 & array_obj_ref_350_word_address_0 & array_obj_ref_338_word_address_0 & array_obj_ref_354_word_address_0 & array_obj_ref_366_word_address_0;
      data_in <= array_obj_ref_342_data_0 & array_obj_ref_326_data_0 & array_obj_ref_330_data_0 & array_obj_ref_318_data_0 & array_obj_ref_358_data_0 & array_obj_ref_362_data_0 & array_obj_ref_334_data_0 & array_obj_ref_346_data_0 & array_obj_ref_310_data_0 & array_obj_ref_314_data_0 & array_obj_ref_322_data_0 & array_obj_ref_350_data_0 & array_obj_ref_338_data_0 & array_obj_ref_354_data_0 & array_obj_ref_366_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 15,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(3 downto 0),
          mdata => memory_space_4_sr_data(7 downto 0),
          mtag => memory_space_4_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr2;
architecture Default of default_initializer_xx_xstr2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr2_CP_1341_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_380_store_0_ack_1 : boolean;
  signal array_obj_ref_372_store_0_req_1 : boolean;
  signal array_obj_ref_408_gather_scatter_req_0 : boolean;
  signal array_obj_ref_420_store_0_req_0 : boolean;
  signal array_obj_ref_424_store_0_req_1 : boolean;
  signal array_obj_ref_412_store_0_req_0 : boolean;
  signal array_obj_ref_412_store_0_ack_0 : boolean;
  signal array_obj_ref_408_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_416_gather_scatter_req_0 : boolean;
  signal array_obj_ref_392_store_0_ack_0 : boolean;
  signal array_obj_ref_388_store_0_req_1 : boolean;
  signal array_obj_ref_416_store_0_req_1 : boolean;
  signal array_obj_ref_412_store_0_req_1 : boolean;
  signal array_obj_ref_376_store_0_req_0 : boolean;
  signal array_obj_ref_424_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_384_store_0_ack_1 : boolean;
  signal array_obj_ref_372_gather_scatter_req_0 : boolean;
  signal array_obj_ref_380_store_0_req_0 : boolean;
  signal array_obj_ref_420_gather_scatter_req_0 : boolean;
  signal array_obj_ref_408_store_0_req_1 : boolean;
  signal array_obj_ref_388_gather_scatter_req_0 : boolean;
  signal array_obj_ref_416_store_0_req_0 : boolean;
  signal array_obj_ref_384_store_0_req_1 : boolean;
  signal array_obj_ref_416_store_0_ack_1 : boolean;
  signal array_obj_ref_392_store_0_req_0 : boolean;
  signal array_obj_ref_372_store_0_req_0 : boolean;
  signal array_obj_ref_380_store_0_ack_0 : boolean;
  signal array_obj_ref_424_store_0_ack_0 : boolean;
  signal array_obj_ref_392_store_0_req_1 : boolean;
  signal array_obj_ref_420_store_0_ack_1 : boolean;
  signal array_obj_ref_416_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_388_store_0_ack_1 : boolean;
  signal array_obj_ref_380_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_380_gather_scatter_req_0 : boolean;
  signal array_obj_ref_408_store_0_ack_1 : boolean;
  signal array_obj_ref_392_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_380_store_0_req_1 : boolean;
  signal array_obj_ref_408_store_0_ack_0 : boolean;
  signal array_obj_ref_376_store_0_ack_1 : boolean;
  signal array_obj_ref_388_store_0_ack_0 : boolean;
  signal array_obj_ref_376_store_0_ack_0 : boolean;
  signal array_obj_ref_424_gather_scatter_req_0 : boolean;
  signal array_obj_ref_384_store_0_req_0 : boolean;
  signal array_obj_ref_376_gather_scatter_req_0 : boolean;
  signal array_obj_ref_388_store_0_req_0 : boolean;
  signal array_obj_ref_416_store_0_ack_0 : boolean;
  signal array_obj_ref_392_gather_scatter_req_0 : boolean;
  signal array_obj_ref_428_gather_scatter_req_0 : boolean;
  signal array_obj_ref_392_store_0_ack_1 : boolean;
  signal array_obj_ref_428_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_408_store_0_req_0 : boolean;
  signal array_obj_ref_412_gather_scatter_req_0 : boolean;
  signal array_obj_ref_420_store_0_req_1 : boolean;
  signal array_obj_ref_372_store_0_ack_0 : boolean;
  signal array_obj_ref_412_store_0_ack_1 : boolean;
  signal array_obj_ref_384_store_0_ack_0 : boolean;
  signal array_obj_ref_372_store_0_ack_1 : boolean;
  signal array_obj_ref_376_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_372_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_420_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_420_store_0_ack_0 : boolean;
  signal array_obj_ref_412_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_424_store_0_req_0 : boolean;
  signal array_obj_ref_376_store_0_req_1 : boolean;
  signal array_obj_ref_404_store_0_ack_1 : boolean;
  signal array_obj_ref_404_store_0_req_1 : boolean;
  signal array_obj_ref_388_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_404_store_0_ack_0 : boolean;
  signal array_obj_ref_404_store_0_req_0 : boolean;
  signal array_obj_ref_404_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_404_gather_scatter_req_0 : boolean;
  signal array_obj_ref_400_store_0_ack_1 : boolean;
  signal array_obj_ref_384_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_400_store_0_req_1 : boolean;
  signal array_obj_ref_400_store_0_ack_0 : boolean;
  signal array_obj_ref_400_store_0_req_0 : boolean;
  signal array_obj_ref_400_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_400_gather_scatter_req_0 : boolean;
  signal array_obj_ref_384_gather_scatter_req_0 : boolean;
  signal array_obj_ref_396_store_0_ack_1 : boolean;
  signal array_obj_ref_396_store_0_req_1 : boolean;
  signal array_obj_ref_396_store_0_ack_0 : boolean;
  signal array_obj_ref_396_store_0_req_0 : boolean;
  signal array_obj_ref_396_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_396_gather_scatter_req_0 : boolean;
  signal array_obj_ref_424_store_0_ack_1 : boolean;
  signal array_obj_ref_428_store_0_ack_1 : boolean;
  signal array_obj_ref_428_store_0_req_1 : boolean;
  signal array_obj_ref_428_store_0_ack_0 : boolean;
  signal array_obj_ref_428_store_0_req_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 15 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr2_CP_1341: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_372_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_372_gather_scatter_ack_0;
    array_obj_ref_372_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_372_store_0_ack_0;
    array_obj_ref_372_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_372_store_0_ack_1;
    array_obj_ref_376_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_376_gather_scatter_ack_0;
    array_obj_ref_376_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_376_store_0_ack_0;
    array_obj_ref_376_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_376_store_0_ack_1;
    array_obj_ref_380_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_380_gather_scatter_ack_0;
    array_obj_ref_380_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_380_store_0_ack_0;
    array_obj_ref_380_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_380_store_0_ack_1;
    array_obj_ref_384_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_384_gather_scatter_ack_0;
    array_obj_ref_384_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_384_store_0_ack_0;
    array_obj_ref_384_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_384_store_0_ack_1;
    array_obj_ref_388_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_388_gather_scatter_ack_0;
    array_obj_ref_388_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_388_store_0_ack_0;
    array_obj_ref_388_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_388_store_0_ack_1;
    array_obj_ref_392_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_392_gather_scatter_ack_0;
    array_obj_ref_392_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_392_store_0_ack_0;
    array_obj_ref_392_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_392_store_0_ack_1;
    array_obj_ref_396_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_396_gather_scatter_ack_0;
    array_obj_ref_396_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_396_store_0_ack_0;
    array_obj_ref_396_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_396_store_0_ack_1;
    array_obj_ref_400_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_400_gather_scatter_ack_0;
    array_obj_ref_400_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_400_store_0_ack_0;
    array_obj_ref_400_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_400_store_0_ack_1;
    array_obj_ref_404_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_404_gather_scatter_ack_0;
    array_obj_ref_404_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_404_store_0_ack_0;
    array_obj_ref_404_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_404_store_0_ack_1;
    array_obj_ref_408_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_408_gather_scatter_ack_0;
    array_obj_ref_408_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_408_store_0_ack_0;
    array_obj_ref_408_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_408_store_0_ack_1;
    array_obj_ref_412_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_412_gather_scatter_ack_0;
    array_obj_ref_412_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_412_store_0_ack_0;
    array_obj_ref_412_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_412_store_0_ack_1;
    array_obj_ref_416_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_416_gather_scatter_ack_0;
    array_obj_ref_416_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_416_store_0_ack_0;
    array_obj_ref_416_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_416_store_0_ack_1;
    array_obj_ref_420_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_420_gather_scatter_ack_0;
    array_obj_ref_420_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_420_store_0_ack_0;
    array_obj_ref_420_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_420_store_0_ack_1;
    array_obj_ref_424_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_424_gather_scatter_ack_0;
    array_obj_ref_424_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_424_store_0_ack_0;
    array_obj_ref_424_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_424_store_0_ack_1;
    array_obj_ref_428_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_428_gather_scatter_ack_0;
    array_obj_ref_428_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_428_store_0_ack_0;
    array_obj_ref_428_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_428_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_372_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_372_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_376_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_376_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_380_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_380_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_384_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_384_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_388_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_388_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_392_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_392_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_396_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_396_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_400_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_400_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_404_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_404_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_408_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_408_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_412_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_412_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_416_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_416_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_420_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_420_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_424_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_424_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_428_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_428_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_373_wire_constant : std_logic_vector(7 downto 0);
    signal expr_377_wire_constant : std_logic_vector(7 downto 0);
    signal expr_381_wire_constant : std_logic_vector(7 downto 0);
    signal expr_385_wire_constant : std_logic_vector(7 downto 0);
    signal expr_389_wire_constant : std_logic_vector(7 downto 0);
    signal expr_393_wire_constant : std_logic_vector(7 downto 0);
    signal expr_397_wire_constant : std_logic_vector(7 downto 0);
    signal expr_401_wire_constant : std_logic_vector(7 downto 0);
    signal expr_405_wire_constant : std_logic_vector(7 downto 0);
    signal expr_409_wire_constant : std_logic_vector(7 downto 0);
    signal expr_413_wire_constant : std_logic_vector(7 downto 0);
    signal expr_417_wire_constant : std_logic_vector(7 downto 0);
    signal expr_421_wire_constant : std_logic_vector(7 downto 0);
    signal expr_425_wire_constant : std_logic_vector(7 downto 0);
    signal expr_429_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_372_word_address_0 <= "0000";
    array_obj_ref_376_word_address_0 <= "0001";
    array_obj_ref_380_word_address_0 <= "0010";
    array_obj_ref_384_word_address_0 <= "0011";
    array_obj_ref_388_word_address_0 <= "0100";
    array_obj_ref_392_word_address_0 <= "0101";
    array_obj_ref_396_word_address_0 <= "0110";
    array_obj_ref_400_word_address_0 <= "0111";
    array_obj_ref_404_word_address_0 <= "1000";
    array_obj_ref_408_word_address_0 <= "1001";
    array_obj_ref_412_word_address_0 <= "1010";
    array_obj_ref_416_word_address_0 <= "1011";
    array_obj_ref_420_word_address_0 <= "1100";
    array_obj_ref_424_word_address_0 <= "1101";
    array_obj_ref_428_word_address_0 <= "1110";
    expr_373_wire_constant <= "01100110";
    expr_377_wire_constant <= "01110010";
    expr_381_wire_constant <= "01100101";
    expr_385_wire_constant <= "01100101";
    expr_389_wire_constant <= "01011111";
    expr_393_wire_constant <= "01110001";
    expr_397_wire_constant <= "01110101";
    expr_401_wire_constant <= "01100101";
    expr_405_wire_constant <= "01110101";
    expr_409_wire_constant <= "01100101";
    expr_413_wire_constant <= "01011111";
    expr_417_wire_constant <= "01100111";
    expr_421_wire_constant <= "01100101";
    expr_425_wire_constant <= "01110100";
    expr_429_wire_constant <= "00000000";
    array_obj_ref_372_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_372_gather_scatter_ack_0 <= array_obj_ref_372_gather_scatter_req_0;
      aggregated_sig <= expr_373_wire_constant;
      array_obj_ref_372_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_376_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_376_gather_scatter_ack_0 <= array_obj_ref_376_gather_scatter_req_0;
      aggregated_sig <= expr_377_wire_constant;
      array_obj_ref_376_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_380_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_380_gather_scatter_ack_0 <= array_obj_ref_380_gather_scatter_req_0;
      aggregated_sig <= expr_381_wire_constant;
      array_obj_ref_380_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_384_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_384_gather_scatter_ack_0 <= array_obj_ref_384_gather_scatter_req_0;
      aggregated_sig <= expr_385_wire_constant;
      array_obj_ref_384_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_388_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_388_gather_scatter_ack_0 <= array_obj_ref_388_gather_scatter_req_0;
      aggregated_sig <= expr_389_wire_constant;
      array_obj_ref_388_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_392_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_392_gather_scatter_ack_0 <= array_obj_ref_392_gather_scatter_req_0;
      aggregated_sig <= expr_393_wire_constant;
      array_obj_ref_392_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_396_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_396_gather_scatter_ack_0 <= array_obj_ref_396_gather_scatter_req_0;
      aggregated_sig <= expr_397_wire_constant;
      array_obj_ref_396_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_400_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_400_gather_scatter_ack_0 <= array_obj_ref_400_gather_scatter_req_0;
      aggregated_sig <= expr_401_wire_constant;
      array_obj_ref_400_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_404_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_404_gather_scatter_ack_0 <= array_obj_ref_404_gather_scatter_req_0;
      aggregated_sig <= expr_405_wire_constant;
      array_obj_ref_404_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_408_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_408_gather_scatter_ack_0 <= array_obj_ref_408_gather_scatter_req_0;
      aggregated_sig <= expr_409_wire_constant;
      array_obj_ref_408_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_412_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_412_gather_scatter_ack_0 <= array_obj_ref_412_gather_scatter_req_0;
      aggregated_sig <= expr_413_wire_constant;
      array_obj_ref_412_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_416_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_416_gather_scatter_ack_0 <= array_obj_ref_416_gather_scatter_req_0;
      aggregated_sig <= expr_417_wire_constant;
      array_obj_ref_416_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_420_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_420_gather_scatter_ack_0 <= array_obj_ref_420_gather_scatter_req_0;
      aggregated_sig <= expr_421_wire_constant;
      array_obj_ref_420_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_424_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_424_gather_scatter_ack_0 <= array_obj_ref_424_gather_scatter_req_0;
      aggregated_sig <= expr_425_wire_constant;
      array_obj_ref_424_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_428_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_428_gather_scatter_ack_0 <= array_obj_ref_428_gather_scatter_req_0;
      aggregated_sig <= expr_429_wire_constant;
      array_obj_ref_428_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_384_store_0 array_obj_ref_388_store_0 array_obj_ref_408_store_0 array_obj_ref_376_store_0 array_obj_ref_424_store_0 array_obj_ref_412_store_0 array_obj_ref_416_store_0 array_obj_ref_404_store_0 array_obj_ref_372_store_0 array_obj_ref_420_store_0 array_obj_ref_396_store_0 array_obj_ref_400_store_0 array_obj_ref_392_store_0 array_obj_ref_428_store_0 array_obj_ref_380_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(59 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_384_store_0_req_0;
      reqL(13) <= array_obj_ref_388_store_0_req_0;
      reqL(12) <= array_obj_ref_408_store_0_req_0;
      reqL(11) <= array_obj_ref_376_store_0_req_0;
      reqL(10) <= array_obj_ref_424_store_0_req_0;
      reqL(9) <= array_obj_ref_412_store_0_req_0;
      reqL(8) <= array_obj_ref_416_store_0_req_0;
      reqL(7) <= array_obj_ref_404_store_0_req_0;
      reqL(6) <= array_obj_ref_372_store_0_req_0;
      reqL(5) <= array_obj_ref_420_store_0_req_0;
      reqL(4) <= array_obj_ref_396_store_0_req_0;
      reqL(3) <= array_obj_ref_400_store_0_req_0;
      reqL(2) <= array_obj_ref_392_store_0_req_0;
      reqL(1) <= array_obj_ref_428_store_0_req_0;
      reqL(0) <= array_obj_ref_380_store_0_req_0;
      array_obj_ref_384_store_0_ack_0 <= ackL(14);
      array_obj_ref_388_store_0_ack_0 <= ackL(13);
      array_obj_ref_408_store_0_ack_0 <= ackL(12);
      array_obj_ref_376_store_0_ack_0 <= ackL(11);
      array_obj_ref_424_store_0_ack_0 <= ackL(10);
      array_obj_ref_412_store_0_ack_0 <= ackL(9);
      array_obj_ref_416_store_0_ack_0 <= ackL(8);
      array_obj_ref_404_store_0_ack_0 <= ackL(7);
      array_obj_ref_372_store_0_ack_0 <= ackL(6);
      array_obj_ref_420_store_0_ack_0 <= ackL(5);
      array_obj_ref_396_store_0_ack_0 <= ackL(4);
      array_obj_ref_400_store_0_ack_0 <= ackL(3);
      array_obj_ref_392_store_0_ack_0 <= ackL(2);
      array_obj_ref_428_store_0_ack_0 <= ackL(1);
      array_obj_ref_380_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_384_store_0_req_1;
      reqR(13) <= array_obj_ref_388_store_0_req_1;
      reqR(12) <= array_obj_ref_408_store_0_req_1;
      reqR(11) <= array_obj_ref_376_store_0_req_1;
      reqR(10) <= array_obj_ref_424_store_0_req_1;
      reqR(9) <= array_obj_ref_412_store_0_req_1;
      reqR(8) <= array_obj_ref_416_store_0_req_1;
      reqR(7) <= array_obj_ref_404_store_0_req_1;
      reqR(6) <= array_obj_ref_372_store_0_req_1;
      reqR(5) <= array_obj_ref_420_store_0_req_1;
      reqR(4) <= array_obj_ref_396_store_0_req_1;
      reqR(3) <= array_obj_ref_400_store_0_req_1;
      reqR(2) <= array_obj_ref_392_store_0_req_1;
      reqR(1) <= array_obj_ref_428_store_0_req_1;
      reqR(0) <= array_obj_ref_380_store_0_req_1;
      array_obj_ref_384_store_0_ack_1 <= ackR(14);
      array_obj_ref_388_store_0_ack_1 <= ackR(13);
      array_obj_ref_408_store_0_ack_1 <= ackR(12);
      array_obj_ref_376_store_0_ack_1 <= ackR(11);
      array_obj_ref_424_store_0_ack_1 <= ackR(10);
      array_obj_ref_412_store_0_ack_1 <= ackR(9);
      array_obj_ref_416_store_0_ack_1 <= ackR(8);
      array_obj_ref_404_store_0_ack_1 <= ackR(7);
      array_obj_ref_372_store_0_ack_1 <= ackR(6);
      array_obj_ref_420_store_0_ack_1 <= ackR(5);
      array_obj_ref_396_store_0_ack_1 <= ackR(4);
      array_obj_ref_400_store_0_ack_1 <= ackR(3);
      array_obj_ref_392_store_0_ack_1 <= ackR(2);
      array_obj_ref_428_store_0_ack_1 <= ackR(1);
      array_obj_ref_380_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_384_word_address_0 & array_obj_ref_388_word_address_0 & array_obj_ref_408_word_address_0 & array_obj_ref_376_word_address_0 & array_obj_ref_424_word_address_0 & array_obj_ref_412_word_address_0 & array_obj_ref_416_word_address_0 & array_obj_ref_404_word_address_0 & array_obj_ref_372_word_address_0 & array_obj_ref_420_word_address_0 & array_obj_ref_396_word_address_0 & array_obj_ref_400_word_address_0 & array_obj_ref_392_word_address_0 & array_obj_ref_428_word_address_0 & array_obj_ref_380_word_address_0;
      data_in <= array_obj_ref_384_data_0 & array_obj_ref_388_data_0 & array_obj_ref_408_data_0 & array_obj_ref_376_data_0 & array_obj_ref_424_data_0 & array_obj_ref_412_data_0 & array_obj_ref_416_data_0 & array_obj_ref_404_data_0 & array_obj_ref_372_data_0 & array_obj_ref_420_data_0 & array_obj_ref_396_data_0 & array_obj_ref_400_data_0 & array_obj_ref_392_data_0 & array_obj_ref_428_data_0 & array_obj_ref_380_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 15,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(3 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr3 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr3;
architecture Default of default_initializer_xx_xstr3 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr3_CP_1659_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_434_gather_scatter_req_0 : boolean;
  signal array_obj_ref_434_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_434_store_0_req_0 : boolean;
  signal array_obj_ref_434_store_0_ack_0 : boolean;
  signal array_obj_ref_434_store_0_req_1 : boolean;
  signal array_obj_ref_434_store_0_ack_1 : boolean;
  signal array_obj_ref_438_gather_scatter_req_0 : boolean;
  signal array_obj_ref_438_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_0 : boolean;
  signal array_obj_ref_438_store_0_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_1 : boolean;
  signal array_obj_ref_438_store_0_ack_1 : boolean;
  signal array_obj_ref_442_gather_scatter_req_0 : boolean;
  signal array_obj_ref_442_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_442_store_0_req_0 : boolean;
  signal array_obj_ref_442_store_0_ack_0 : boolean;
  signal array_obj_ref_442_store_0_req_1 : boolean;
  signal array_obj_ref_442_store_0_ack_1 : boolean;
  signal array_obj_ref_446_gather_scatter_req_0 : boolean;
  signal array_obj_ref_446_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_446_store_0_req_0 : boolean;
  signal array_obj_ref_446_store_0_ack_0 : boolean;
  signal array_obj_ref_446_store_0_req_1 : boolean;
  signal array_obj_ref_446_store_0_ack_1 : boolean;
  signal array_obj_ref_450_gather_scatter_req_0 : boolean;
  signal array_obj_ref_450_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_450_store_0_req_0 : boolean;
  signal array_obj_ref_450_store_0_ack_0 : boolean;
  signal array_obj_ref_450_store_0_req_1 : boolean;
  signal array_obj_ref_450_store_0_ack_1 : boolean;
  signal array_obj_ref_454_gather_scatter_req_0 : boolean;
  signal array_obj_ref_454_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_454_store_0_req_0 : boolean;
  signal array_obj_ref_454_store_0_ack_0 : boolean;
  signal array_obj_ref_454_store_0_req_1 : boolean;
  signal array_obj_ref_454_store_0_ack_1 : boolean;
  signal array_obj_ref_458_gather_scatter_req_0 : boolean;
  signal array_obj_ref_458_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_0 : boolean;
  signal array_obj_ref_458_store_0_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_1 : boolean;
  signal array_obj_ref_458_store_0_ack_1 : boolean;
  signal array_obj_ref_462_gather_scatter_req_0 : boolean;
  signal array_obj_ref_462_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_462_store_0_req_0 : boolean;
  signal array_obj_ref_462_store_0_ack_0 : boolean;
  signal array_obj_ref_462_store_0_req_1 : boolean;
  signal array_obj_ref_462_store_0_ack_1 : boolean;
  signal array_obj_ref_466_gather_scatter_req_0 : boolean;
  signal array_obj_ref_466_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_466_store_0_req_0 : boolean;
  signal array_obj_ref_466_store_0_ack_0 : boolean;
  signal array_obj_ref_466_store_0_req_1 : boolean;
  signal array_obj_ref_466_store_0_ack_1 : boolean;
  signal array_obj_ref_470_gather_scatter_req_0 : boolean;
  signal array_obj_ref_470_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_470_store_0_req_0 : boolean;
  signal array_obj_ref_470_store_0_ack_0 : boolean;
  signal array_obj_ref_470_store_0_req_1 : boolean;
  signal array_obj_ref_470_store_0_ack_1 : boolean;
  signal array_obj_ref_474_gather_scatter_req_0 : boolean;
  signal array_obj_ref_474_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_474_store_0_req_0 : boolean;
  signal array_obj_ref_474_store_0_ack_0 : boolean;
  signal array_obj_ref_474_store_0_req_1 : boolean;
  signal array_obj_ref_474_store_0_ack_1 : boolean;
  signal array_obj_ref_478_gather_scatter_req_0 : boolean;
  signal array_obj_ref_478_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_478_store_0_req_0 : boolean;
  signal array_obj_ref_478_store_0_ack_0 : boolean;
  signal array_obj_ref_478_store_0_req_1 : boolean;
  signal array_obj_ref_478_store_0_ack_1 : boolean;
  signal array_obj_ref_482_gather_scatter_req_0 : boolean;
  signal array_obj_ref_482_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_482_store_0_req_0 : boolean;
  signal array_obj_ref_482_store_0_ack_0 : boolean;
  signal array_obj_ref_482_store_0_req_1 : boolean;
  signal array_obj_ref_482_store_0_ack_1 : boolean;
  signal array_obj_ref_486_gather_scatter_req_0 : boolean;
  signal array_obj_ref_486_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_486_store_0_req_0 : boolean;
  signal array_obj_ref_486_store_0_ack_0 : boolean;
  signal array_obj_ref_486_store_0_req_1 : boolean;
  signal array_obj_ref_486_store_0_ack_1 : boolean;
  signal array_obj_ref_490_gather_scatter_req_0 : boolean;
  signal array_obj_ref_490_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_490_store_0_req_0 : boolean;
  signal array_obj_ref_490_store_0_ack_0 : boolean;
  signal array_obj_ref_490_store_0_req_1 : boolean;
  signal array_obj_ref_490_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 15 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr3_CP_1659: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_434_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_434_gather_scatter_ack_0;
    array_obj_ref_434_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_434_store_0_ack_0;
    array_obj_ref_434_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_434_store_0_ack_1;
    array_obj_ref_438_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_438_gather_scatter_ack_0;
    array_obj_ref_438_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_438_store_0_ack_0;
    array_obj_ref_438_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_438_store_0_ack_1;
    array_obj_ref_442_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_442_gather_scatter_ack_0;
    array_obj_ref_442_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_442_store_0_ack_0;
    array_obj_ref_442_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_442_store_0_ack_1;
    array_obj_ref_446_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_446_gather_scatter_ack_0;
    array_obj_ref_446_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_446_store_0_ack_0;
    array_obj_ref_446_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_446_store_0_ack_1;
    array_obj_ref_450_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_450_gather_scatter_ack_0;
    array_obj_ref_450_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_450_store_0_ack_0;
    array_obj_ref_450_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_450_store_0_ack_1;
    array_obj_ref_454_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_454_gather_scatter_ack_0;
    array_obj_ref_454_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_454_store_0_ack_0;
    array_obj_ref_454_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_454_store_0_ack_1;
    array_obj_ref_458_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_458_gather_scatter_ack_0;
    array_obj_ref_458_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_458_store_0_ack_0;
    array_obj_ref_458_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_458_store_0_ack_1;
    array_obj_ref_462_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_462_gather_scatter_ack_0;
    array_obj_ref_462_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_462_store_0_ack_0;
    array_obj_ref_462_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_462_store_0_ack_1;
    array_obj_ref_466_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_466_gather_scatter_ack_0;
    array_obj_ref_466_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_466_store_0_ack_0;
    array_obj_ref_466_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_466_store_0_ack_1;
    array_obj_ref_470_gather_scatter_req_0 <= cp_elements(27);
    cp_elements(28) <= array_obj_ref_470_gather_scatter_ack_0;
    array_obj_ref_470_store_0_req_0 <= cp_elements(28);
    cp_elements(29) <= array_obj_ref_470_store_0_ack_0;
    array_obj_ref_470_store_0_req_1 <= cp_elements(29);
    cp_elements(30) <= array_obj_ref_470_store_0_ack_1;
    array_obj_ref_474_gather_scatter_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_474_gather_scatter_ack_0;
    array_obj_ref_474_store_0_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_474_store_0_ack_0;
    array_obj_ref_474_store_0_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_474_store_0_ack_1;
    array_obj_ref_478_gather_scatter_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_478_gather_scatter_ack_0;
    array_obj_ref_478_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_478_store_0_ack_0;
    array_obj_ref_478_store_0_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_478_store_0_ack_1;
    array_obj_ref_482_gather_scatter_req_0 <= cp_elements(36);
    cp_elements(37) <= array_obj_ref_482_gather_scatter_ack_0;
    array_obj_ref_482_store_0_req_0 <= cp_elements(37);
    cp_elements(38) <= array_obj_ref_482_store_0_ack_0;
    array_obj_ref_482_store_0_req_1 <= cp_elements(38);
    cp_elements(39) <= array_obj_ref_482_store_0_ack_1;
    array_obj_ref_486_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= array_obj_ref_486_gather_scatter_ack_0;
    array_obj_ref_486_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= array_obj_ref_486_store_0_ack_0;
    array_obj_ref_486_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= array_obj_ref_486_store_0_ack_1;
    array_obj_ref_490_gather_scatter_req_0 <= cp_elements(42);
    cp_elements(43) <= array_obj_ref_490_gather_scatter_ack_0;
    array_obj_ref_490_store_0_req_0 <= cp_elements(43);
    cp_elements(44) <= array_obj_ref_490_store_0_ack_0;
    array_obj_ref_490_store_0_req_1 <= cp_elements(44);
    cp_elements(45) <= array_obj_ref_490_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_434_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_434_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_438_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_438_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_442_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_442_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_446_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_446_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_450_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_450_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_454_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_454_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_458_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_458_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_462_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_462_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_466_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_466_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_470_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_470_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_474_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_474_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_478_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_478_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_482_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_482_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_486_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_486_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_490_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_490_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_435_wire_constant : std_logic_vector(7 downto 0);
    signal expr_439_wire_constant : std_logic_vector(7 downto 0);
    signal expr_443_wire_constant : std_logic_vector(7 downto 0);
    signal expr_447_wire_constant : std_logic_vector(7 downto 0);
    signal expr_451_wire_constant : std_logic_vector(7 downto 0);
    signal expr_455_wire_constant : std_logic_vector(7 downto 0);
    signal expr_459_wire_constant : std_logic_vector(7 downto 0);
    signal expr_463_wire_constant : std_logic_vector(7 downto 0);
    signal expr_467_wire_constant : std_logic_vector(7 downto 0);
    signal expr_471_wire_constant : std_logic_vector(7 downto 0);
    signal expr_475_wire_constant : std_logic_vector(7 downto 0);
    signal expr_479_wire_constant : std_logic_vector(7 downto 0);
    signal expr_483_wire_constant : std_logic_vector(7 downto 0);
    signal expr_487_wire_constant : std_logic_vector(7 downto 0);
    signal expr_491_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_434_word_address_0 <= "0000";
    array_obj_ref_438_word_address_0 <= "0001";
    array_obj_ref_442_word_address_0 <= "0010";
    array_obj_ref_446_word_address_0 <= "0011";
    array_obj_ref_450_word_address_0 <= "0100";
    array_obj_ref_454_word_address_0 <= "0101";
    array_obj_ref_458_word_address_0 <= "0110";
    array_obj_ref_462_word_address_0 <= "0111";
    array_obj_ref_466_word_address_0 <= "1000";
    array_obj_ref_470_word_address_0 <= "1001";
    array_obj_ref_474_word_address_0 <= "1010";
    array_obj_ref_478_word_address_0 <= "1011";
    array_obj_ref_482_word_address_0 <= "1100";
    array_obj_ref_486_word_address_0 <= "1101";
    array_obj_ref_490_word_address_0 <= "1110";
    expr_435_wire_constant <= "01100110";
    expr_439_wire_constant <= "01110010";
    expr_443_wire_constant <= "01100101";
    expr_447_wire_constant <= "01100101";
    expr_451_wire_constant <= "01011111";
    expr_455_wire_constant <= "01110001";
    expr_459_wire_constant <= "01110101";
    expr_463_wire_constant <= "01100101";
    expr_467_wire_constant <= "01110101";
    expr_471_wire_constant <= "01100101";
    expr_475_wire_constant <= "01011111";
    expr_479_wire_constant <= "01110000";
    expr_483_wire_constant <= "01110101";
    expr_487_wire_constant <= "01110100";
    expr_491_wire_constant <= "00000000";
    array_obj_ref_434_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_434_gather_scatter_ack_0 <= array_obj_ref_434_gather_scatter_req_0;
      aggregated_sig <= expr_435_wire_constant;
      array_obj_ref_434_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_438_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_438_gather_scatter_ack_0 <= array_obj_ref_438_gather_scatter_req_0;
      aggregated_sig <= expr_439_wire_constant;
      array_obj_ref_438_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_442_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_442_gather_scatter_ack_0 <= array_obj_ref_442_gather_scatter_req_0;
      aggregated_sig <= expr_443_wire_constant;
      array_obj_ref_442_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_446_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_446_gather_scatter_ack_0 <= array_obj_ref_446_gather_scatter_req_0;
      aggregated_sig <= expr_447_wire_constant;
      array_obj_ref_446_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_450_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_450_gather_scatter_ack_0 <= array_obj_ref_450_gather_scatter_req_0;
      aggregated_sig <= expr_451_wire_constant;
      array_obj_ref_450_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_454_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_454_gather_scatter_ack_0 <= array_obj_ref_454_gather_scatter_req_0;
      aggregated_sig <= expr_455_wire_constant;
      array_obj_ref_454_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_458_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_458_gather_scatter_ack_0 <= array_obj_ref_458_gather_scatter_req_0;
      aggregated_sig <= expr_459_wire_constant;
      array_obj_ref_458_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_462_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_462_gather_scatter_ack_0 <= array_obj_ref_462_gather_scatter_req_0;
      aggregated_sig <= expr_463_wire_constant;
      array_obj_ref_462_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_466_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_466_gather_scatter_ack_0 <= array_obj_ref_466_gather_scatter_req_0;
      aggregated_sig <= expr_467_wire_constant;
      array_obj_ref_466_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_470_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_470_gather_scatter_ack_0 <= array_obj_ref_470_gather_scatter_req_0;
      aggregated_sig <= expr_471_wire_constant;
      array_obj_ref_470_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_474_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_474_gather_scatter_ack_0 <= array_obj_ref_474_gather_scatter_req_0;
      aggregated_sig <= expr_475_wire_constant;
      array_obj_ref_474_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_478_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_478_gather_scatter_ack_0 <= array_obj_ref_478_gather_scatter_req_0;
      aggregated_sig <= expr_479_wire_constant;
      array_obj_ref_478_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_482_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_482_gather_scatter_ack_0 <= array_obj_ref_482_gather_scatter_req_0;
      aggregated_sig <= expr_483_wire_constant;
      array_obj_ref_482_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_486_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_486_gather_scatter_ack_0 <= array_obj_ref_486_gather_scatter_req_0;
      aggregated_sig <= expr_487_wire_constant;
      array_obj_ref_486_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_490_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_490_gather_scatter_ack_0 <= array_obj_ref_490_gather_scatter_req_0;
      aggregated_sig <= expr_491_wire_constant;
      array_obj_ref_490_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_458_store_0 array_obj_ref_490_store_0 array_obj_ref_486_store_0 array_obj_ref_478_store_0 array_obj_ref_482_store_0 array_obj_ref_438_store_0 array_obj_ref_434_store_0 array_obj_ref_470_store_0 array_obj_ref_462_store_0 array_obj_ref_442_store_0 array_obj_ref_466_store_0 array_obj_ref_474_store_0 array_obj_ref_454_store_0 array_obj_ref_450_store_0 array_obj_ref_446_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(59 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_458_store_0_req_0;
      reqL(13) <= array_obj_ref_490_store_0_req_0;
      reqL(12) <= array_obj_ref_486_store_0_req_0;
      reqL(11) <= array_obj_ref_478_store_0_req_0;
      reqL(10) <= array_obj_ref_482_store_0_req_0;
      reqL(9) <= array_obj_ref_438_store_0_req_0;
      reqL(8) <= array_obj_ref_434_store_0_req_0;
      reqL(7) <= array_obj_ref_470_store_0_req_0;
      reqL(6) <= array_obj_ref_462_store_0_req_0;
      reqL(5) <= array_obj_ref_442_store_0_req_0;
      reqL(4) <= array_obj_ref_466_store_0_req_0;
      reqL(3) <= array_obj_ref_474_store_0_req_0;
      reqL(2) <= array_obj_ref_454_store_0_req_0;
      reqL(1) <= array_obj_ref_450_store_0_req_0;
      reqL(0) <= array_obj_ref_446_store_0_req_0;
      array_obj_ref_458_store_0_ack_0 <= ackL(14);
      array_obj_ref_490_store_0_ack_0 <= ackL(13);
      array_obj_ref_486_store_0_ack_0 <= ackL(12);
      array_obj_ref_478_store_0_ack_0 <= ackL(11);
      array_obj_ref_482_store_0_ack_0 <= ackL(10);
      array_obj_ref_438_store_0_ack_0 <= ackL(9);
      array_obj_ref_434_store_0_ack_0 <= ackL(8);
      array_obj_ref_470_store_0_ack_0 <= ackL(7);
      array_obj_ref_462_store_0_ack_0 <= ackL(6);
      array_obj_ref_442_store_0_ack_0 <= ackL(5);
      array_obj_ref_466_store_0_ack_0 <= ackL(4);
      array_obj_ref_474_store_0_ack_0 <= ackL(3);
      array_obj_ref_454_store_0_ack_0 <= ackL(2);
      array_obj_ref_450_store_0_ack_0 <= ackL(1);
      array_obj_ref_446_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_458_store_0_req_1;
      reqR(13) <= array_obj_ref_490_store_0_req_1;
      reqR(12) <= array_obj_ref_486_store_0_req_1;
      reqR(11) <= array_obj_ref_478_store_0_req_1;
      reqR(10) <= array_obj_ref_482_store_0_req_1;
      reqR(9) <= array_obj_ref_438_store_0_req_1;
      reqR(8) <= array_obj_ref_434_store_0_req_1;
      reqR(7) <= array_obj_ref_470_store_0_req_1;
      reqR(6) <= array_obj_ref_462_store_0_req_1;
      reqR(5) <= array_obj_ref_442_store_0_req_1;
      reqR(4) <= array_obj_ref_466_store_0_req_1;
      reqR(3) <= array_obj_ref_474_store_0_req_1;
      reqR(2) <= array_obj_ref_454_store_0_req_1;
      reqR(1) <= array_obj_ref_450_store_0_req_1;
      reqR(0) <= array_obj_ref_446_store_0_req_1;
      array_obj_ref_458_store_0_ack_1 <= ackR(14);
      array_obj_ref_490_store_0_ack_1 <= ackR(13);
      array_obj_ref_486_store_0_ack_1 <= ackR(12);
      array_obj_ref_478_store_0_ack_1 <= ackR(11);
      array_obj_ref_482_store_0_ack_1 <= ackR(10);
      array_obj_ref_438_store_0_ack_1 <= ackR(9);
      array_obj_ref_434_store_0_ack_1 <= ackR(8);
      array_obj_ref_470_store_0_ack_1 <= ackR(7);
      array_obj_ref_462_store_0_ack_1 <= ackR(6);
      array_obj_ref_442_store_0_ack_1 <= ackR(5);
      array_obj_ref_466_store_0_ack_1 <= ackR(4);
      array_obj_ref_474_store_0_ack_1 <= ackR(3);
      array_obj_ref_454_store_0_ack_1 <= ackR(2);
      array_obj_ref_450_store_0_ack_1 <= ackR(1);
      array_obj_ref_446_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_458_word_address_0 & array_obj_ref_490_word_address_0 & array_obj_ref_486_word_address_0 & array_obj_ref_478_word_address_0 & array_obj_ref_482_word_address_0 & array_obj_ref_438_word_address_0 & array_obj_ref_434_word_address_0 & array_obj_ref_470_word_address_0 & array_obj_ref_462_word_address_0 & array_obj_ref_442_word_address_0 & array_obj_ref_466_word_address_0 & array_obj_ref_474_word_address_0 & array_obj_ref_454_word_address_0 & array_obj_ref_450_word_address_0 & array_obj_ref_446_word_address_0;
      data_in <= array_obj_ref_458_data_0 & array_obj_ref_490_data_0 & array_obj_ref_486_data_0 & array_obj_ref_478_data_0 & array_obj_ref_482_data_0 & array_obj_ref_438_data_0 & array_obj_ref_434_data_0 & array_obj_ref_470_data_0 & array_obj_ref_462_data_0 & array_obj_ref_442_data_0 & array_obj_ref_466_data_0 & array_obj_ref_474_data_0 & array_obj_ref_454_data_0 & array_obj_ref_450_data_0 & array_obj_ref_446_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 15,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(3 downto 0),
          mdata => memory_space_6_sr_data(7 downto 0),
          mtag => memory_space_6_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr4;
architecture Default of default_initializer_xx_xstr4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr4_CP_1977_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_516_store_0_ack_0 : boolean;
  signal array_obj_ref_504_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_516_gather_scatter_req_0 : boolean;
  signal array_obj_ref_524_store_0_req_1 : boolean;
  signal array_obj_ref_524_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_516_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_520_gather_scatter_req_0 : boolean;
  signal array_obj_ref_520_store_0_req_0 : boolean;
  signal array_obj_ref_508_store_0_req_1 : boolean;
  signal array_obj_ref_508_store_0_ack_1 : boolean;
  signal array_obj_ref_504_gather_scatter_req_0 : boolean;
  signal array_obj_ref_508_store_0_ack_0 : boolean;
  signal array_obj_ref_500_gather_scatter_req_0 : boolean;
  signal array_obj_ref_524_store_0_ack_0 : boolean;
  signal array_obj_ref_520_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_512_store_0_req_1 : boolean;
  signal array_obj_ref_500_store_0_ack_0 : boolean;
  signal array_obj_ref_508_store_0_req_0 : boolean;
  signal array_obj_ref_520_store_0_ack_0 : boolean;
  signal array_obj_ref_500_store_0_ack_1 : boolean;
  signal array_obj_ref_516_store_0_req_0 : boolean;
  signal array_obj_ref_500_store_0_req_1 : boolean;
  signal array_obj_ref_500_store_0_req_0 : boolean;
  signal array_obj_ref_524_gather_scatter_req_0 : boolean;
  signal array_obj_ref_504_store_0_req_0 : boolean;
  signal array_obj_ref_516_store_0_ack_1 : boolean;
  signal array_obj_ref_504_store_0_ack_0 : boolean;
  signal array_obj_ref_504_store_0_req_1 : boolean;
  signal array_obj_ref_504_store_0_ack_1 : boolean;
  signal array_obj_ref_512_gather_scatter_req_0 : boolean;
  signal array_obj_ref_512_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_500_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_516_store_0_req_1 : boolean;
  signal array_obj_ref_512_store_0_req_0 : boolean;
  signal array_obj_ref_508_gather_scatter_req_0 : boolean;
  signal array_obj_ref_512_store_0_ack_1 : boolean;
  signal array_obj_ref_508_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_512_store_0_ack_0 : boolean;
  signal array_obj_ref_496_store_0_ack_1 : boolean;
  signal array_obj_ref_496_store_0_req_1 : boolean;
  signal array_obj_ref_524_store_0_ack_1 : boolean;
  signal array_obj_ref_496_store_0_ack_0 : boolean;
  signal array_obj_ref_496_store_0_req_0 : boolean;
  signal array_obj_ref_524_store_0_req_0 : boolean;
  signal array_obj_ref_496_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_496_gather_scatter_req_0 : boolean;
  signal array_obj_ref_520_store_0_ack_1 : boolean;
  signal array_obj_ref_520_store_0_req_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 8 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr4_CP_1977: Block -- control-path 
    signal cp_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(24);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(24), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_496_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_496_gather_scatter_ack_0;
    array_obj_ref_496_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_496_store_0_ack_0;
    array_obj_ref_496_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_496_store_0_ack_1;
    array_obj_ref_500_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_500_gather_scatter_ack_0;
    array_obj_ref_500_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_500_store_0_ack_0;
    array_obj_ref_500_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_500_store_0_ack_1;
    array_obj_ref_504_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_504_gather_scatter_ack_0;
    array_obj_ref_504_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_504_store_0_ack_0;
    array_obj_ref_504_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_504_store_0_ack_1;
    array_obj_ref_508_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_508_gather_scatter_ack_0;
    array_obj_ref_508_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_508_store_0_ack_0;
    array_obj_ref_508_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_508_store_0_ack_1;
    array_obj_ref_512_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_512_gather_scatter_ack_0;
    array_obj_ref_512_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_512_store_0_ack_0;
    array_obj_ref_512_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_512_store_0_ack_1;
    array_obj_ref_516_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_516_gather_scatter_ack_0;
    array_obj_ref_516_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_516_store_0_ack_0;
    array_obj_ref_516_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_516_store_0_ack_1;
    array_obj_ref_520_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_520_gather_scatter_ack_0;
    array_obj_ref_520_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_520_store_0_ack_0;
    array_obj_ref_520_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_520_store_0_ack_1;
    array_obj_ref_524_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_524_gather_scatter_ack_0;
    array_obj_ref_524_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_524_store_0_ack_0;
    array_obj_ref_524_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_524_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_496_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_496_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_500_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_500_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_504_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_504_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_508_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_508_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_512_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_512_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_516_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_516_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_520_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_520_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_524_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_524_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_497_wire_constant : std_logic_vector(7 downto 0);
    signal expr_501_wire_constant : std_logic_vector(7 downto 0);
    signal expr_505_wire_constant : std_logic_vector(7 downto 0);
    signal expr_509_wire_constant : std_logic_vector(7 downto 0);
    signal expr_513_wire_constant : std_logic_vector(7 downto 0);
    signal expr_517_wire_constant : std_logic_vector(7 downto 0);
    signal expr_521_wire_constant : std_logic_vector(7 downto 0);
    signal expr_525_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_496_word_address_0 <= "0000";
    array_obj_ref_500_word_address_0 <= "0001";
    array_obj_ref_504_word_address_0 <= "0010";
    array_obj_ref_508_word_address_0 <= "0011";
    array_obj_ref_512_word_address_0 <= "0100";
    array_obj_ref_516_word_address_0 <= "0101";
    array_obj_ref_520_word_address_0 <= "0110";
    array_obj_ref_524_word_address_0 <= "0111";
    expr_497_wire_constant <= "01101001";
    expr_501_wire_constant <= "01101110";
    expr_505_wire_constant <= "01011111";
    expr_509_wire_constant <= "01100100";
    expr_513_wire_constant <= "01100001";
    expr_517_wire_constant <= "01110100";
    expr_521_wire_constant <= "01100001";
    expr_525_wire_constant <= "00000000";
    array_obj_ref_496_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_496_gather_scatter_ack_0 <= array_obj_ref_496_gather_scatter_req_0;
      aggregated_sig <= expr_497_wire_constant;
      array_obj_ref_496_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_500_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_500_gather_scatter_ack_0 <= array_obj_ref_500_gather_scatter_req_0;
      aggregated_sig <= expr_501_wire_constant;
      array_obj_ref_500_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_504_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_504_gather_scatter_ack_0 <= array_obj_ref_504_gather_scatter_req_0;
      aggregated_sig <= expr_505_wire_constant;
      array_obj_ref_504_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_508_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_508_gather_scatter_ack_0 <= array_obj_ref_508_gather_scatter_req_0;
      aggregated_sig <= expr_509_wire_constant;
      array_obj_ref_508_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_512_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_512_gather_scatter_ack_0 <= array_obj_ref_512_gather_scatter_req_0;
      aggregated_sig <= expr_513_wire_constant;
      array_obj_ref_512_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_516_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_516_gather_scatter_ack_0 <= array_obj_ref_516_gather_scatter_req_0;
      aggregated_sig <= expr_517_wire_constant;
      array_obj_ref_516_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_520_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_520_gather_scatter_ack_0 <= array_obj_ref_520_gather_scatter_req_0;
      aggregated_sig <= expr_521_wire_constant;
      array_obj_ref_520_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_524_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_524_gather_scatter_ack_0 <= array_obj_ref_524_gather_scatter_req_0;
      aggregated_sig <= expr_525_wire_constant;
      array_obj_ref_524_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_524_store_0 array_obj_ref_496_store_0 array_obj_ref_508_store_0 array_obj_ref_516_store_0 array_obj_ref_504_store_0 array_obj_ref_500_store_0 array_obj_ref_512_store_0 array_obj_ref_520_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(31 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= array_obj_ref_524_store_0_req_0;
      reqL(6) <= array_obj_ref_496_store_0_req_0;
      reqL(5) <= array_obj_ref_508_store_0_req_0;
      reqL(4) <= array_obj_ref_516_store_0_req_0;
      reqL(3) <= array_obj_ref_504_store_0_req_0;
      reqL(2) <= array_obj_ref_500_store_0_req_0;
      reqL(1) <= array_obj_ref_512_store_0_req_0;
      reqL(0) <= array_obj_ref_520_store_0_req_0;
      array_obj_ref_524_store_0_ack_0 <= ackL(7);
      array_obj_ref_496_store_0_ack_0 <= ackL(6);
      array_obj_ref_508_store_0_ack_0 <= ackL(5);
      array_obj_ref_516_store_0_ack_0 <= ackL(4);
      array_obj_ref_504_store_0_ack_0 <= ackL(3);
      array_obj_ref_500_store_0_ack_0 <= ackL(2);
      array_obj_ref_512_store_0_ack_0 <= ackL(1);
      array_obj_ref_520_store_0_ack_0 <= ackL(0);
      reqR(7) <= array_obj_ref_524_store_0_req_1;
      reqR(6) <= array_obj_ref_496_store_0_req_1;
      reqR(5) <= array_obj_ref_508_store_0_req_1;
      reqR(4) <= array_obj_ref_516_store_0_req_1;
      reqR(3) <= array_obj_ref_504_store_0_req_1;
      reqR(2) <= array_obj_ref_500_store_0_req_1;
      reqR(1) <= array_obj_ref_512_store_0_req_1;
      reqR(0) <= array_obj_ref_520_store_0_req_1;
      array_obj_ref_524_store_0_ack_1 <= ackR(7);
      array_obj_ref_496_store_0_ack_1 <= ackR(6);
      array_obj_ref_508_store_0_ack_1 <= ackR(5);
      array_obj_ref_516_store_0_ack_1 <= ackR(4);
      array_obj_ref_504_store_0_ack_1 <= ackR(3);
      array_obj_ref_500_store_0_ack_1 <= ackR(2);
      array_obj_ref_512_store_0_ack_1 <= ackR(1);
      array_obj_ref_520_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_524_word_address_0 & array_obj_ref_496_word_address_0 & array_obj_ref_508_word_address_0 & array_obj_ref_516_word_address_0 & array_obj_ref_504_word_address_0 & array_obj_ref_500_word_address_0 & array_obj_ref_512_word_address_0 & array_obj_ref_520_word_address_0;
      data_in <= array_obj_ref_524_data_0 & array_obj_ref_496_data_0 & array_obj_ref_508_data_0 & array_obj_ref_516_data_0 & array_obj_ref_504_data_0 & array_obj_ref_500_data_0 & array_obj_ref_512_data_0 & array_obj_ref_520_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(3 downto 0),
          mdata => memory_space_7_sr_data(7 downto 0),
          mtag => memory_space_7_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr5 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr5;
architecture Default of default_initializer_xx_xstr5 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr5_CP_2148_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_542_store_0_req_0 : boolean;
  signal array_obj_ref_542_store_0_ack_0 : boolean;
  signal array_obj_ref_542_store_0_req_1 : boolean;
  signal array_obj_ref_542_gather_scatter_req_0 : boolean;
  signal array_obj_ref_542_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_538_gather_scatter_req_0 : boolean;
  signal array_obj_ref_538_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_538_store_0_req_0 : boolean;
  signal array_obj_ref_530_gather_scatter_req_0 : boolean;
  signal array_obj_ref_538_store_0_ack_0 : boolean;
  signal array_obj_ref_538_store_0_req_1 : boolean;
  signal array_obj_ref_538_store_0_ack_1 : boolean;
  signal array_obj_ref_554_gather_scatter_req_0 : boolean;
  signal array_obj_ref_554_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_534_store_0_req_1 : boolean;
  signal array_obj_ref_534_store_0_ack_1 : boolean;
  signal array_obj_ref_550_store_0_req_0 : boolean;
  signal array_obj_ref_550_store_0_ack_0 : boolean;
  signal array_obj_ref_550_store_0_req_1 : boolean;
  signal array_obj_ref_550_store_0_ack_1 : boolean;
  signal array_obj_ref_534_store_0_req_0 : boolean;
  signal array_obj_ref_534_store_0_ack_0 : boolean;
  signal array_obj_ref_550_gather_scatter_req_0 : boolean;
  signal array_obj_ref_550_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_534_gather_scatter_req_0 : boolean;
  signal array_obj_ref_534_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_546_store_0_ack_0 : boolean;
  signal array_obj_ref_546_store_0_req_1 : boolean;
  signal array_obj_ref_546_store_0_ack_1 : boolean;
  signal array_obj_ref_546_gather_scatter_req_0 : boolean;
  signal array_obj_ref_546_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_546_store_0_req_0 : boolean;
  signal array_obj_ref_530_store_0_ack_1 : boolean;
  signal array_obj_ref_542_store_0_ack_1 : boolean;
  signal array_obj_ref_530_store_0_req_0 : boolean;
  signal array_obj_ref_530_store_0_ack_0 : boolean;
  signal array_obj_ref_530_store_0_req_1 : boolean;
  signal array_obj_ref_554_store_0_req_0 : boolean;
  signal array_obj_ref_554_store_0_ack_0 : boolean;
  signal array_obj_ref_554_store_0_req_1 : boolean;
  signal array_obj_ref_554_store_0_ack_1 : boolean;
  signal array_obj_ref_530_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_558_gather_scatter_req_0 : boolean;
  signal array_obj_ref_558_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_558_store_0_req_0 : boolean;
  signal array_obj_ref_558_store_0_ack_0 : boolean;
  signal array_obj_ref_558_store_0_req_1 : boolean;
  signal array_obj_ref_558_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 8 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr5_CP_2148: Block -- control-path 
    signal cp_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(24);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(24), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_530_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_530_gather_scatter_ack_0;
    array_obj_ref_530_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_530_store_0_ack_0;
    array_obj_ref_530_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_530_store_0_ack_1;
    array_obj_ref_534_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_534_gather_scatter_ack_0;
    array_obj_ref_534_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_534_store_0_ack_0;
    array_obj_ref_534_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_534_store_0_ack_1;
    array_obj_ref_538_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_538_gather_scatter_ack_0;
    array_obj_ref_538_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_538_store_0_ack_0;
    array_obj_ref_538_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_538_store_0_ack_1;
    array_obj_ref_542_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_542_gather_scatter_ack_0;
    array_obj_ref_542_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_542_store_0_ack_0;
    array_obj_ref_542_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_542_store_0_ack_1;
    array_obj_ref_546_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_546_gather_scatter_ack_0;
    array_obj_ref_546_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_546_store_0_ack_0;
    array_obj_ref_546_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_546_store_0_ack_1;
    array_obj_ref_550_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_550_gather_scatter_ack_0;
    array_obj_ref_550_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_550_store_0_ack_0;
    array_obj_ref_550_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_550_store_0_ack_1;
    array_obj_ref_554_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_554_gather_scatter_ack_0;
    array_obj_ref_554_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_554_store_0_ack_0;
    array_obj_ref_554_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_554_store_0_ack_1;
    array_obj_ref_558_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_558_gather_scatter_ack_0;
    array_obj_ref_558_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_558_store_0_ack_0;
    array_obj_ref_558_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_558_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_530_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_530_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_534_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_534_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_538_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_538_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_542_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_542_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_546_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_546_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_550_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_550_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_554_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_554_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_558_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_558_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_531_wire_constant : std_logic_vector(7 downto 0);
    signal expr_535_wire_constant : std_logic_vector(7 downto 0);
    signal expr_539_wire_constant : std_logic_vector(7 downto 0);
    signal expr_543_wire_constant : std_logic_vector(7 downto 0);
    signal expr_547_wire_constant : std_logic_vector(7 downto 0);
    signal expr_551_wire_constant : std_logic_vector(7 downto 0);
    signal expr_555_wire_constant : std_logic_vector(7 downto 0);
    signal expr_559_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_530_word_address_0 <= "0000";
    array_obj_ref_534_word_address_0 <= "0001";
    array_obj_ref_538_word_address_0 <= "0010";
    array_obj_ref_542_word_address_0 <= "0011";
    array_obj_ref_546_word_address_0 <= "0100";
    array_obj_ref_550_word_address_0 <= "0101";
    array_obj_ref_554_word_address_0 <= "0110";
    array_obj_ref_558_word_address_0 <= "0111";
    expr_531_wire_constant <= "01101001";
    expr_535_wire_constant <= "01101110";
    expr_539_wire_constant <= "01011111";
    expr_543_wire_constant <= "01100011";
    expr_547_wire_constant <= "01110100";
    expr_551_wire_constant <= "01110010";
    expr_555_wire_constant <= "01101100";
    expr_559_wire_constant <= "00000000";
    array_obj_ref_530_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_530_gather_scatter_ack_0 <= array_obj_ref_530_gather_scatter_req_0;
      aggregated_sig <= expr_531_wire_constant;
      array_obj_ref_530_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_534_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_534_gather_scatter_ack_0 <= array_obj_ref_534_gather_scatter_req_0;
      aggregated_sig <= expr_535_wire_constant;
      array_obj_ref_534_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_538_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_538_gather_scatter_ack_0 <= array_obj_ref_538_gather_scatter_req_0;
      aggregated_sig <= expr_539_wire_constant;
      array_obj_ref_538_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_542_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_542_gather_scatter_ack_0 <= array_obj_ref_542_gather_scatter_req_0;
      aggregated_sig <= expr_543_wire_constant;
      array_obj_ref_542_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_546_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_546_gather_scatter_ack_0 <= array_obj_ref_546_gather_scatter_req_0;
      aggregated_sig <= expr_547_wire_constant;
      array_obj_ref_546_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_550_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_550_gather_scatter_ack_0 <= array_obj_ref_550_gather_scatter_req_0;
      aggregated_sig <= expr_551_wire_constant;
      array_obj_ref_550_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_554_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_554_gather_scatter_ack_0 <= array_obj_ref_554_gather_scatter_req_0;
      aggregated_sig <= expr_555_wire_constant;
      array_obj_ref_554_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_558_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_558_gather_scatter_ack_0 <= array_obj_ref_558_gather_scatter_req_0;
      aggregated_sig <= expr_559_wire_constant;
      array_obj_ref_558_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_530_store_0 array_obj_ref_534_store_0 array_obj_ref_538_store_0 array_obj_ref_542_store_0 array_obj_ref_546_store_0 array_obj_ref_550_store_0 array_obj_ref_554_store_0 array_obj_ref_558_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(31 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= array_obj_ref_530_store_0_req_0;
      reqL(6) <= array_obj_ref_534_store_0_req_0;
      reqL(5) <= array_obj_ref_538_store_0_req_0;
      reqL(4) <= array_obj_ref_542_store_0_req_0;
      reqL(3) <= array_obj_ref_546_store_0_req_0;
      reqL(2) <= array_obj_ref_550_store_0_req_0;
      reqL(1) <= array_obj_ref_554_store_0_req_0;
      reqL(0) <= array_obj_ref_558_store_0_req_0;
      array_obj_ref_530_store_0_ack_0 <= ackL(7);
      array_obj_ref_534_store_0_ack_0 <= ackL(6);
      array_obj_ref_538_store_0_ack_0 <= ackL(5);
      array_obj_ref_542_store_0_ack_0 <= ackL(4);
      array_obj_ref_546_store_0_ack_0 <= ackL(3);
      array_obj_ref_550_store_0_ack_0 <= ackL(2);
      array_obj_ref_554_store_0_ack_0 <= ackL(1);
      array_obj_ref_558_store_0_ack_0 <= ackL(0);
      reqR(7) <= array_obj_ref_530_store_0_req_1;
      reqR(6) <= array_obj_ref_534_store_0_req_1;
      reqR(5) <= array_obj_ref_538_store_0_req_1;
      reqR(4) <= array_obj_ref_542_store_0_req_1;
      reqR(3) <= array_obj_ref_546_store_0_req_1;
      reqR(2) <= array_obj_ref_550_store_0_req_1;
      reqR(1) <= array_obj_ref_554_store_0_req_1;
      reqR(0) <= array_obj_ref_558_store_0_req_1;
      array_obj_ref_530_store_0_ack_1 <= ackR(7);
      array_obj_ref_534_store_0_ack_1 <= ackR(6);
      array_obj_ref_538_store_0_ack_1 <= ackR(5);
      array_obj_ref_542_store_0_ack_1 <= ackR(4);
      array_obj_ref_546_store_0_ack_1 <= ackR(3);
      array_obj_ref_550_store_0_ack_1 <= ackR(2);
      array_obj_ref_554_store_0_ack_1 <= ackR(1);
      array_obj_ref_558_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_530_word_address_0 & array_obj_ref_534_word_address_0 & array_obj_ref_538_word_address_0 & array_obj_ref_542_word_address_0 & array_obj_ref_546_word_address_0 & array_obj_ref_550_word_address_0 & array_obj_ref_554_word_address_0 & array_obj_ref_558_word_address_0;
      data_in <= array_obj_ref_530_data_0 & array_obj_ref_534_data_0 & array_obj_ref_538_data_0 & array_obj_ref_542_data_0 & array_obj_ref_546_data_0 & array_obj_ref_550_data_0 & array_obj_ref_554_data_0 & array_obj_ref_558_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(3 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr6 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_9_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_9_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_9_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr6;
architecture Default of default_initializer_xx_xstr6 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr6_CP_2319_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_564_gather_scatter_req_0 : boolean;
  signal array_obj_ref_564_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_564_store_0_req_0 : boolean;
  signal array_obj_ref_564_store_0_ack_0 : boolean;
  signal array_obj_ref_564_store_0_req_1 : boolean;
  signal array_obj_ref_564_store_0_ack_1 : boolean;
  signal array_obj_ref_568_gather_scatter_req_0 : boolean;
  signal array_obj_ref_568_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_568_store_0_req_0 : boolean;
  signal array_obj_ref_568_store_0_ack_0 : boolean;
  signal array_obj_ref_568_store_0_req_1 : boolean;
  signal array_obj_ref_568_store_0_ack_1 : boolean;
  signal array_obj_ref_572_gather_scatter_req_0 : boolean;
  signal array_obj_ref_572_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_572_store_0_req_0 : boolean;
  signal array_obj_ref_572_store_0_ack_0 : boolean;
  signal array_obj_ref_572_store_0_req_1 : boolean;
  signal array_obj_ref_572_store_0_ack_1 : boolean;
  signal array_obj_ref_576_gather_scatter_req_0 : boolean;
  signal array_obj_ref_576_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_576_store_0_req_0 : boolean;
  signal array_obj_ref_576_store_0_ack_0 : boolean;
  signal array_obj_ref_576_store_0_req_1 : boolean;
  signal array_obj_ref_576_store_0_ack_1 : boolean;
  signal array_obj_ref_580_gather_scatter_req_0 : boolean;
  signal array_obj_ref_580_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_580_store_0_req_0 : boolean;
  signal array_obj_ref_580_store_0_ack_0 : boolean;
  signal array_obj_ref_580_store_0_req_1 : boolean;
  signal array_obj_ref_580_store_0_ack_1 : boolean;
  signal array_obj_ref_584_gather_scatter_req_0 : boolean;
  signal array_obj_ref_584_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_584_store_0_req_0 : boolean;
  signal array_obj_ref_584_store_0_ack_0 : boolean;
  signal array_obj_ref_584_store_0_req_1 : boolean;
  signal array_obj_ref_584_store_0_ack_1 : boolean;
  signal array_obj_ref_588_gather_scatter_req_0 : boolean;
  signal array_obj_ref_588_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_588_store_0_req_0 : boolean;
  signal array_obj_ref_588_store_0_ack_0 : boolean;
  signal array_obj_ref_588_store_0_req_1 : boolean;
  signal array_obj_ref_588_store_0_ack_1 : boolean;
  signal array_obj_ref_592_gather_scatter_req_0 : boolean;
  signal array_obj_ref_592_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_592_store_0_req_0 : boolean;
  signal array_obj_ref_592_store_0_ack_0 : boolean;
  signal array_obj_ref_592_store_0_req_1 : boolean;
  signal array_obj_ref_592_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 8 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr6_CP_2319: Block -- control-path 
    signal cp_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(24);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(24), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_564_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_564_gather_scatter_ack_0;
    array_obj_ref_564_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_564_store_0_ack_0;
    array_obj_ref_564_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_564_store_0_ack_1;
    array_obj_ref_568_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_568_gather_scatter_ack_0;
    array_obj_ref_568_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_568_store_0_ack_0;
    array_obj_ref_568_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_568_store_0_ack_1;
    array_obj_ref_572_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_572_gather_scatter_ack_0;
    array_obj_ref_572_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_572_store_0_ack_0;
    array_obj_ref_572_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_572_store_0_ack_1;
    array_obj_ref_576_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_576_gather_scatter_ack_0;
    array_obj_ref_576_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_576_store_0_ack_0;
    array_obj_ref_576_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_576_store_0_ack_1;
    array_obj_ref_580_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_580_gather_scatter_ack_0;
    array_obj_ref_580_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_580_store_0_ack_0;
    array_obj_ref_580_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_580_store_0_ack_1;
    array_obj_ref_584_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_584_gather_scatter_ack_0;
    array_obj_ref_584_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_584_store_0_ack_0;
    array_obj_ref_584_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_584_store_0_ack_1;
    array_obj_ref_588_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_588_gather_scatter_ack_0;
    array_obj_ref_588_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_588_store_0_ack_0;
    array_obj_ref_588_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_588_store_0_ack_1;
    array_obj_ref_592_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_592_gather_scatter_ack_0;
    array_obj_ref_592_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_592_store_0_ack_0;
    array_obj_ref_592_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_592_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_564_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_564_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_568_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_568_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_572_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_572_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_576_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_576_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_580_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_580_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_584_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_584_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_588_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_588_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_592_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_592_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_565_wire_constant : std_logic_vector(7 downto 0);
    signal expr_569_wire_constant : std_logic_vector(7 downto 0);
    signal expr_573_wire_constant : std_logic_vector(7 downto 0);
    signal expr_577_wire_constant : std_logic_vector(7 downto 0);
    signal expr_581_wire_constant : std_logic_vector(7 downto 0);
    signal expr_585_wire_constant : std_logic_vector(7 downto 0);
    signal expr_589_wire_constant : std_logic_vector(7 downto 0);
    signal expr_593_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_564_word_address_0 <= "0000";
    array_obj_ref_568_word_address_0 <= "0001";
    array_obj_ref_572_word_address_0 <= "0010";
    array_obj_ref_576_word_address_0 <= "0011";
    array_obj_ref_580_word_address_0 <= "0100";
    array_obj_ref_584_word_address_0 <= "0101";
    array_obj_ref_588_word_address_0 <= "0110";
    array_obj_ref_592_word_address_0 <= "0111";
    expr_565_wire_constant <= "01101101";
    expr_569_wire_constant <= "01101001";
    expr_573_wire_constant <= "01100100";
    expr_577_wire_constant <= "01110000";
    expr_581_wire_constant <= "01101001";
    expr_585_wire_constant <= "01110000";
    expr_589_wire_constant <= "01100101";
    expr_593_wire_constant <= "00000000";
    array_obj_ref_564_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_564_gather_scatter_ack_0 <= array_obj_ref_564_gather_scatter_req_0;
      aggregated_sig <= expr_565_wire_constant;
      array_obj_ref_564_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_568_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_568_gather_scatter_ack_0 <= array_obj_ref_568_gather_scatter_req_0;
      aggregated_sig <= expr_569_wire_constant;
      array_obj_ref_568_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_572_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_572_gather_scatter_ack_0 <= array_obj_ref_572_gather_scatter_req_0;
      aggregated_sig <= expr_573_wire_constant;
      array_obj_ref_572_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_576_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_576_gather_scatter_ack_0 <= array_obj_ref_576_gather_scatter_req_0;
      aggregated_sig <= expr_577_wire_constant;
      array_obj_ref_576_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_580_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_580_gather_scatter_ack_0 <= array_obj_ref_580_gather_scatter_req_0;
      aggregated_sig <= expr_581_wire_constant;
      array_obj_ref_580_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_584_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_584_gather_scatter_ack_0 <= array_obj_ref_584_gather_scatter_req_0;
      aggregated_sig <= expr_585_wire_constant;
      array_obj_ref_584_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_588_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_588_gather_scatter_ack_0 <= array_obj_ref_588_gather_scatter_req_0;
      aggregated_sig <= expr_589_wire_constant;
      array_obj_ref_588_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_592_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_592_gather_scatter_ack_0 <= array_obj_ref_592_gather_scatter_req_0;
      aggregated_sig <= expr_593_wire_constant;
      array_obj_ref_592_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_580_store_0 array_obj_ref_592_store_0 array_obj_ref_588_store_0 array_obj_ref_568_store_0 array_obj_ref_572_store_0 array_obj_ref_576_store_0 array_obj_ref_564_store_0 array_obj_ref_584_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(31 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= array_obj_ref_580_store_0_req_0;
      reqL(6) <= array_obj_ref_592_store_0_req_0;
      reqL(5) <= array_obj_ref_588_store_0_req_0;
      reqL(4) <= array_obj_ref_568_store_0_req_0;
      reqL(3) <= array_obj_ref_572_store_0_req_0;
      reqL(2) <= array_obj_ref_576_store_0_req_0;
      reqL(1) <= array_obj_ref_564_store_0_req_0;
      reqL(0) <= array_obj_ref_584_store_0_req_0;
      array_obj_ref_580_store_0_ack_0 <= ackL(7);
      array_obj_ref_592_store_0_ack_0 <= ackL(6);
      array_obj_ref_588_store_0_ack_0 <= ackL(5);
      array_obj_ref_568_store_0_ack_0 <= ackL(4);
      array_obj_ref_572_store_0_ack_0 <= ackL(3);
      array_obj_ref_576_store_0_ack_0 <= ackL(2);
      array_obj_ref_564_store_0_ack_0 <= ackL(1);
      array_obj_ref_584_store_0_ack_0 <= ackL(0);
      reqR(7) <= array_obj_ref_580_store_0_req_1;
      reqR(6) <= array_obj_ref_592_store_0_req_1;
      reqR(5) <= array_obj_ref_588_store_0_req_1;
      reqR(4) <= array_obj_ref_568_store_0_req_1;
      reqR(3) <= array_obj_ref_572_store_0_req_1;
      reqR(2) <= array_obj_ref_576_store_0_req_1;
      reqR(1) <= array_obj_ref_564_store_0_req_1;
      reqR(0) <= array_obj_ref_584_store_0_req_1;
      array_obj_ref_580_store_0_ack_1 <= ackR(7);
      array_obj_ref_592_store_0_ack_1 <= ackR(6);
      array_obj_ref_588_store_0_ack_1 <= ackR(5);
      array_obj_ref_568_store_0_ack_1 <= ackR(4);
      array_obj_ref_572_store_0_ack_1 <= ackR(3);
      array_obj_ref_576_store_0_ack_1 <= ackR(2);
      array_obj_ref_564_store_0_ack_1 <= ackR(1);
      array_obj_ref_584_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_580_word_address_0 & array_obj_ref_592_word_address_0 & array_obj_ref_588_word_address_0 & array_obj_ref_568_word_address_0 & array_obj_ref_572_word_address_0 & array_obj_ref_576_word_address_0 & array_obj_ref_564_word_address_0 & array_obj_ref_584_word_address_0;
      data_in <= array_obj_ref_580_data_0 & array_obj_ref_592_data_0 & array_obj_ref_588_data_0 & array_obj_ref_568_data_0 & array_obj_ref_572_data_0 & array_obj_ref_576_data_0 & array_obj_ref_564_data_0 & array_obj_ref_584_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(3 downto 0),
          mdata => memory_space_9_sr_data(7 downto 0),
          mtag => memory_space_9_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr7 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_10_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_10_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_10_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr7;
architecture Default of default_initializer_xx_xstr7 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr7_CP_2490_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_618_store_0_req_1 : boolean;
  signal array_obj_ref_622_store_0_req_1 : boolean;
  signal array_obj_ref_618_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_618_store_0_req_0 : boolean;
  signal array_obj_ref_602_store_0_req_1 : boolean;
  signal array_obj_ref_622_gather_scatter_req_0 : boolean;
  signal array_obj_ref_606_store_0_req_0 : boolean;
  signal array_obj_ref_606_store_0_ack_0 : boolean;
  signal array_obj_ref_618_store_0_ack_1 : boolean;
  signal array_obj_ref_630_store_0_req_0 : boolean;
  signal array_obj_ref_618_store_0_ack_0 : boolean;
  signal array_obj_ref_610_store_0_req_1 : boolean;
  signal array_obj_ref_610_gather_scatter_req_0 : boolean;
  signal array_obj_ref_622_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_606_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_630_store_0_req_1 : boolean;
  signal array_obj_ref_602_gather_scatter_req_0 : boolean;
  signal array_obj_ref_598_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_614_gather_scatter_req_0 : boolean;
  signal array_obj_ref_626_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_606_store_0_req_1 : boolean;
  signal array_obj_ref_602_store_0_ack_1 : boolean;
  signal array_obj_ref_610_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_626_store_0_req_1 : boolean;
  signal array_obj_ref_606_gather_scatter_req_0 : boolean;
  signal array_obj_ref_622_store_0_req_0 : boolean;
  signal array_obj_ref_622_store_0_ack_1 : boolean;
  signal array_obj_ref_610_store_0_ack_0 : boolean;
  signal array_obj_ref_602_store_0_req_0 : boolean;
  signal array_obj_ref_598_gather_scatter_req_0 : boolean;
  signal array_obj_ref_606_store_0_ack_1 : boolean;
  signal array_obj_ref_610_store_0_req_0 : boolean;
  signal array_obj_ref_610_store_0_ack_1 : boolean;
  signal array_obj_ref_626_gather_scatter_req_0 : boolean;
  signal array_obj_ref_598_store_0_req_1 : boolean;
  signal array_obj_ref_626_store_0_ack_1 : boolean;
  signal array_obj_ref_602_store_0_ack_0 : boolean;
  signal array_obj_ref_618_gather_scatter_req_0 : boolean;
  signal array_obj_ref_622_store_0_ack_0 : boolean;
  signal array_obj_ref_630_store_0_ack_0 : boolean;
  signal array_obj_ref_598_store_0_ack_0 : boolean;
  signal array_obj_ref_626_store_0_req_0 : boolean;
  signal array_obj_ref_598_store_0_req_0 : boolean;
  signal array_obj_ref_598_store_0_ack_1 : boolean;
  signal array_obj_ref_614_store_0_ack_1 : boolean;
  signal array_obj_ref_630_store_0_ack_1 : boolean;
  signal array_obj_ref_626_store_0_ack_0 : boolean;
  signal array_obj_ref_602_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_614_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_630_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_614_store_0_req_0 : boolean;
  signal array_obj_ref_614_store_0_ack_0 : boolean;
  signal array_obj_ref_630_gather_scatter_req_0 : boolean;
  signal array_obj_ref_614_store_0_req_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 9 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr7_CP_2490: Block -- control-path 
    signal cp_elements: BooleanArray(27 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(27);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(27), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_598_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_598_gather_scatter_ack_0;
    array_obj_ref_598_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_598_store_0_ack_0;
    array_obj_ref_598_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_598_store_0_ack_1;
    array_obj_ref_602_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_602_gather_scatter_ack_0;
    array_obj_ref_602_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_602_store_0_ack_0;
    array_obj_ref_602_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_602_store_0_ack_1;
    array_obj_ref_606_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_606_gather_scatter_ack_0;
    array_obj_ref_606_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_606_store_0_ack_0;
    array_obj_ref_606_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_606_store_0_ack_1;
    array_obj_ref_610_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_610_gather_scatter_ack_0;
    array_obj_ref_610_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_610_store_0_ack_0;
    array_obj_ref_610_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_610_store_0_ack_1;
    array_obj_ref_614_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_614_gather_scatter_ack_0;
    array_obj_ref_614_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_614_store_0_ack_0;
    array_obj_ref_614_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_614_store_0_ack_1;
    array_obj_ref_618_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_618_gather_scatter_ack_0;
    array_obj_ref_618_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_618_store_0_ack_0;
    array_obj_ref_618_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_618_store_0_ack_1;
    array_obj_ref_622_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_622_gather_scatter_ack_0;
    array_obj_ref_622_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_622_store_0_ack_0;
    array_obj_ref_622_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_622_store_0_ack_1;
    array_obj_ref_626_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_626_gather_scatter_ack_0;
    array_obj_ref_626_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_626_store_0_ack_0;
    array_obj_ref_626_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_626_store_0_ack_1;
    array_obj_ref_630_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_630_gather_scatter_ack_0;
    array_obj_ref_630_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_630_store_0_ack_0;
    array_obj_ref_630_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_630_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_598_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_598_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_602_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_602_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_606_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_606_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_610_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_610_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_614_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_614_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_618_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_618_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_622_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_622_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_626_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_626_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_630_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_630_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_599_wire_constant : std_logic_vector(7 downto 0);
    signal expr_603_wire_constant : std_logic_vector(7 downto 0);
    signal expr_607_wire_constant : std_logic_vector(7 downto 0);
    signal expr_611_wire_constant : std_logic_vector(7 downto 0);
    signal expr_615_wire_constant : std_logic_vector(7 downto 0);
    signal expr_619_wire_constant : std_logic_vector(7 downto 0);
    signal expr_623_wire_constant : std_logic_vector(7 downto 0);
    signal expr_627_wire_constant : std_logic_vector(7 downto 0);
    signal expr_631_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_598_word_address_0 <= "0000";
    array_obj_ref_602_word_address_0 <= "0001";
    array_obj_ref_606_word_address_0 <= "0010";
    array_obj_ref_610_word_address_0 <= "0011";
    array_obj_ref_614_word_address_0 <= "0100";
    array_obj_ref_618_word_address_0 <= "0101";
    array_obj_ref_622_word_address_0 <= "0110";
    array_obj_ref_626_word_address_0 <= "0111";
    array_obj_ref_630_word_address_0 <= "1000";
    expr_599_wire_constant <= "01101111";
    expr_603_wire_constant <= "01110101";
    expr_607_wire_constant <= "01110100";
    expr_611_wire_constant <= "01011111";
    expr_615_wire_constant <= "01100011";
    expr_619_wire_constant <= "01110100";
    expr_623_wire_constant <= "01110010";
    expr_627_wire_constant <= "01101100";
    expr_631_wire_constant <= "00000000";
    array_obj_ref_598_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_598_gather_scatter_ack_0 <= array_obj_ref_598_gather_scatter_req_0;
      aggregated_sig <= expr_599_wire_constant;
      array_obj_ref_598_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_602_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_602_gather_scatter_ack_0 <= array_obj_ref_602_gather_scatter_req_0;
      aggregated_sig <= expr_603_wire_constant;
      array_obj_ref_602_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_606_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_606_gather_scatter_ack_0 <= array_obj_ref_606_gather_scatter_req_0;
      aggregated_sig <= expr_607_wire_constant;
      array_obj_ref_606_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_610_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_610_gather_scatter_ack_0 <= array_obj_ref_610_gather_scatter_req_0;
      aggregated_sig <= expr_611_wire_constant;
      array_obj_ref_610_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_614_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_614_gather_scatter_ack_0 <= array_obj_ref_614_gather_scatter_req_0;
      aggregated_sig <= expr_615_wire_constant;
      array_obj_ref_614_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_618_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_618_gather_scatter_ack_0 <= array_obj_ref_618_gather_scatter_req_0;
      aggregated_sig <= expr_619_wire_constant;
      array_obj_ref_618_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_622_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_622_gather_scatter_ack_0 <= array_obj_ref_622_gather_scatter_req_0;
      aggregated_sig <= expr_623_wire_constant;
      array_obj_ref_622_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_626_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_626_gather_scatter_ack_0 <= array_obj_ref_626_gather_scatter_req_0;
      aggregated_sig <= expr_627_wire_constant;
      array_obj_ref_626_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_630_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_630_gather_scatter_ack_0 <= array_obj_ref_630_gather_scatter_req_0;
      aggregated_sig <= expr_631_wire_constant;
      array_obj_ref_630_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_602_store_0 array_obj_ref_606_store_0 array_obj_ref_598_store_0 array_obj_ref_618_store_0 array_obj_ref_614_store_0 array_obj_ref_630_store_0 array_obj_ref_626_store_0 array_obj_ref_610_store_0 array_obj_ref_622_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(35 downto 0);
      signal data_in: std_logic_vector(71 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 8 downto 0);
      -- 
    begin -- 
      reqL(8) <= array_obj_ref_602_store_0_req_0;
      reqL(7) <= array_obj_ref_606_store_0_req_0;
      reqL(6) <= array_obj_ref_598_store_0_req_0;
      reqL(5) <= array_obj_ref_618_store_0_req_0;
      reqL(4) <= array_obj_ref_614_store_0_req_0;
      reqL(3) <= array_obj_ref_630_store_0_req_0;
      reqL(2) <= array_obj_ref_626_store_0_req_0;
      reqL(1) <= array_obj_ref_610_store_0_req_0;
      reqL(0) <= array_obj_ref_622_store_0_req_0;
      array_obj_ref_602_store_0_ack_0 <= ackL(8);
      array_obj_ref_606_store_0_ack_0 <= ackL(7);
      array_obj_ref_598_store_0_ack_0 <= ackL(6);
      array_obj_ref_618_store_0_ack_0 <= ackL(5);
      array_obj_ref_614_store_0_ack_0 <= ackL(4);
      array_obj_ref_630_store_0_ack_0 <= ackL(3);
      array_obj_ref_626_store_0_ack_0 <= ackL(2);
      array_obj_ref_610_store_0_ack_0 <= ackL(1);
      array_obj_ref_622_store_0_ack_0 <= ackL(0);
      reqR(8) <= array_obj_ref_602_store_0_req_1;
      reqR(7) <= array_obj_ref_606_store_0_req_1;
      reqR(6) <= array_obj_ref_598_store_0_req_1;
      reqR(5) <= array_obj_ref_618_store_0_req_1;
      reqR(4) <= array_obj_ref_614_store_0_req_1;
      reqR(3) <= array_obj_ref_630_store_0_req_1;
      reqR(2) <= array_obj_ref_626_store_0_req_1;
      reqR(1) <= array_obj_ref_610_store_0_req_1;
      reqR(0) <= array_obj_ref_622_store_0_req_1;
      array_obj_ref_602_store_0_ack_1 <= ackR(8);
      array_obj_ref_606_store_0_ack_1 <= ackR(7);
      array_obj_ref_598_store_0_ack_1 <= ackR(6);
      array_obj_ref_618_store_0_ack_1 <= ackR(5);
      array_obj_ref_614_store_0_ack_1 <= ackR(4);
      array_obj_ref_630_store_0_ack_1 <= ackR(3);
      array_obj_ref_626_store_0_ack_1 <= ackR(2);
      array_obj_ref_610_store_0_ack_1 <= ackR(1);
      array_obj_ref_622_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_602_word_address_0 & array_obj_ref_606_word_address_0 & array_obj_ref_598_word_address_0 & array_obj_ref_618_word_address_0 & array_obj_ref_614_word_address_0 & array_obj_ref_630_word_address_0 & array_obj_ref_626_word_address_0 & array_obj_ref_610_word_address_0 & array_obj_ref_622_word_address_0;
      data_in <= array_obj_ref_602_data_0 & array_obj_ref_606_data_0 & array_obj_ref_598_data_0 & array_obj_ref_618_data_0 & array_obj_ref_614_data_0 & array_obj_ref_630_data_0 & array_obj_ref_626_data_0 & array_obj_ref_610_data_0 & array_obj_ref_622_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 9,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_10_sr_req(0),
          mack => memory_space_10_sr_ack(0),
          maddr => memory_space_10_sr_addr(3 downto 0),
          mdata => memory_space_10_sr_data(7 downto 0),
          mtag => memory_space_10_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 9,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_10_sc_req(0),
          mack => memory_space_10_sc_ack(0),
          mtag => memory_space_10_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity default_initializer_xx_xstr8 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_11_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_11_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_11_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_11_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_11_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_11_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_11_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity default_initializer_xx_xstr8;
architecture Default of default_initializer_xx_xstr8 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal default_initializer_xx_xstr8_CP_2682_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_636_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_640_store_0_ack_1 : boolean;
  signal array_obj_ref_656_store_0_req_1 : boolean;
  signal array_obj_ref_656_store_0_ack_1 : boolean;
  signal array_obj_ref_640_store_0_req_0 : boolean;
  signal array_obj_ref_652_store_0_req_0 : boolean;
  signal array_obj_ref_652_store_0_req_1 : boolean;
  signal array_obj_ref_652_store_0_ack_0 : boolean;
  signal array_obj_ref_640_store_0_req_1 : boolean;
  signal array_obj_ref_640_store_0_ack_0 : boolean;
  signal array_obj_ref_636_gather_scatter_req_0 : boolean;
  signal array_obj_ref_648_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_648_store_0_req_0 : boolean;
  signal array_obj_ref_648_store_0_ack_0 : boolean;
  signal array_obj_ref_636_store_0_ack_1 : boolean;
  signal array_obj_ref_644_store_0_req_1 : boolean;
  signal array_obj_ref_644_store_0_ack_1 : boolean;
  signal array_obj_ref_660_gather_scatter_req_0 : boolean;
  signal array_obj_ref_648_gather_scatter_req_0 : boolean;
  signal array_obj_ref_644_gather_scatter_req_0 : boolean;
  signal array_obj_ref_668_store_0_req_1 : boolean;
  signal array_obj_ref_668_store_0_ack_1 : boolean;
  signal array_obj_ref_648_store_0_req_1 : boolean;
  signal array_obj_ref_664_store_0_ack_1 : boolean;
  signal array_obj_ref_664_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_636_store_0_req_0 : boolean;
  signal array_obj_ref_636_store_0_req_1 : boolean;
  signal array_obj_ref_664_store_0_ack_0 : boolean;
  signal array_obj_ref_664_store_0_req_1 : boolean;
  signal array_obj_ref_664_store_0_req_0 : boolean;
  signal array_obj_ref_664_gather_scatter_req_0 : boolean;
  signal array_obj_ref_668_store_0_req_0 : boolean;
  signal array_obj_ref_668_store_0_ack_0 : boolean;
  signal array_obj_ref_656_store_0_ack_0 : boolean;
  signal array_obj_ref_656_store_0_req_0 : boolean;
  signal array_obj_ref_636_store_0_ack_0 : boolean;
  signal array_obj_ref_660_store_0_ack_1 : boolean;
  signal array_obj_ref_640_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_660_store_0_req_1 : boolean;
  signal array_obj_ref_640_gather_scatter_req_0 : boolean;
  signal array_obj_ref_660_store_0_req_0 : boolean;
  signal array_obj_ref_660_store_0_ack_0 : boolean;
  signal array_obj_ref_660_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_644_store_0_ack_0 : boolean;
  signal array_obj_ref_644_store_0_req_0 : boolean;
  signal array_obj_ref_644_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_652_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_656_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_652_gather_scatter_req_0 : boolean;
  signal array_obj_ref_656_gather_scatter_req_0 : boolean;
  signal array_obj_ref_648_store_0_ack_1 : boolean;
  signal array_obj_ref_652_store_0_ack_1 : boolean;
  signal array_obj_ref_668_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_668_gather_scatter_req_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 9 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  default_initializer_xx_xstr8_CP_2682: Block -- control-path 
    signal cp_elements: BooleanArray(27 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(27);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(27), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    array_obj_ref_636_gather_scatter_req_0 <= cp_elements(0);
    cp_elements(1) <= array_obj_ref_636_gather_scatter_ack_0;
    array_obj_ref_636_store_0_req_0 <= cp_elements(1);
    cp_elements(2) <= array_obj_ref_636_store_0_ack_0;
    array_obj_ref_636_store_0_req_1 <= cp_elements(2);
    cp_elements(3) <= array_obj_ref_636_store_0_ack_1;
    array_obj_ref_640_gather_scatter_req_0 <= cp_elements(3);
    cp_elements(4) <= array_obj_ref_640_gather_scatter_ack_0;
    array_obj_ref_640_store_0_req_0 <= cp_elements(4);
    cp_elements(5) <= array_obj_ref_640_store_0_ack_0;
    array_obj_ref_640_store_0_req_1 <= cp_elements(5);
    cp_elements(6) <= array_obj_ref_640_store_0_ack_1;
    array_obj_ref_644_gather_scatter_req_0 <= cp_elements(6);
    cp_elements(7) <= array_obj_ref_644_gather_scatter_ack_0;
    array_obj_ref_644_store_0_req_0 <= cp_elements(7);
    cp_elements(8) <= array_obj_ref_644_store_0_ack_0;
    array_obj_ref_644_store_0_req_1 <= cp_elements(8);
    cp_elements(9) <= array_obj_ref_644_store_0_ack_1;
    array_obj_ref_648_gather_scatter_req_0 <= cp_elements(9);
    cp_elements(10) <= array_obj_ref_648_gather_scatter_ack_0;
    array_obj_ref_648_store_0_req_0 <= cp_elements(10);
    cp_elements(11) <= array_obj_ref_648_store_0_ack_0;
    array_obj_ref_648_store_0_req_1 <= cp_elements(11);
    cp_elements(12) <= array_obj_ref_648_store_0_ack_1;
    array_obj_ref_652_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_652_gather_scatter_ack_0;
    array_obj_ref_652_store_0_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_652_store_0_ack_0;
    array_obj_ref_652_store_0_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_652_store_0_ack_1;
    array_obj_ref_656_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_656_gather_scatter_ack_0;
    array_obj_ref_656_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_656_store_0_ack_0;
    array_obj_ref_656_store_0_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_656_store_0_ack_1;
    array_obj_ref_660_gather_scatter_req_0 <= cp_elements(18);
    cp_elements(19) <= array_obj_ref_660_gather_scatter_ack_0;
    array_obj_ref_660_store_0_req_0 <= cp_elements(19);
    cp_elements(20) <= array_obj_ref_660_store_0_ack_0;
    array_obj_ref_660_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= array_obj_ref_660_store_0_ack_1;
    array_obj_ref_664_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= array_obj_ref_664_gather_scatter_ack_0;
    array_obj_ref_664_store_0_req_0 <= cp_elements(22);
    cp_elements(23) <= array_obj_ref_664_store_0_ack_0;
    array_obj_ref_664_store_0_req_1 <= cp_elements(23);
    cp_elements(24) <= array_obj_ref_664_store_0_ack_1;
    array_obj_ref_668_gather_scatter_req_0 <= cp_elements(24);
    cp_elements(25) <= array_obj_ref_668_gather_scatter_ack_0;
    array_obj_ref_668_store_0_req_0 <= cp_elements(25);
    cp_elements(26) <= array_obj_ref_668_store_0_ack_0;
    array_obj_ref_668_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= array_obj_ref_668_store_0_ack_1;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_636_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_636_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_640_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_640_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_644_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_644_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_648_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_648_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_652_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_652_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_656_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_656_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_660_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_660_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_664_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_664_word_address_0 : std_logic_vector(3 downto 0);
    signal array_obj_ref_668_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_668_word_address_0 : std_logic_vector(3 downto 0);
    signal expr_637_wire_constant : std_logic_vector(7 downto 0);
    signal expr_641_wire_constant : std_logic_vector(7 downto 0);
    signal expr_645_wire_constant : std_logic_vector(7 downto 0);
    signal expr_649_wire_constant : std_logic_vector(7 downto 0);
    signal expr_653_wire_constant : std_logic_vector(7 downto 0);
    signal expr_657_wire_constant : std_logic_vector(7 downto 0);
    signal expr_661_wire_constant : std_logic_vector(7 downto 0);
    signal expr_665_wire_constant : std_logic_vector(7 downto 0);
    signal expr_669_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_636_word_address_0 <= "0000";
    array_obj_ref_640_word_address_0 <= "0001";
    array_obj_ref_644_word_address_0 <= "0010";
    array_obj_ref_648_word_address_0 <= "0011";
    array_obj_ref_652_word_address_0 <= "0100";
    array_obj_ref_656_word_address_0 <= "0101";
    array_obj_ref_660_word_address_0 <= "0110";
    array_obj_ref_664_word_address_0 <= "0111";
    array_obj_ref_668_word_address_0 <= "1000";
    expr_637_wire_constant <= "01101111";
    expr_641_wire_constant <= "01110101";
    expr_645_wire_constant <= "01110100";
    expr_649_wire_constant <= "01011111";
    expr_653_wire_constant <= "01100100";
    expr_657_wire_constant <= "01100001";
    expr_661_wire_constant <= "01110100";
    expr_665_wire_constant <= "01100001";
    expr_669_wire_constant <= "00000000";
    array_obj_ref_636_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_636_gather_scatter_ack_0 <= array_obj_ref_636_gather_scatter_req_0;
      aggregated_sig <= expr_637_wire_constant;
      array_obj_ref_636_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_640_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_640_gather_scatter_ack_0 <= array_obj_ref_640_gather_scatter_req_0;
      aggregated_sig <= expr_641_wire_constant;
      array_obj_ref_640_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_644_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_644_gather_scatter_ack_0 <= array_obj_ref_644_gather_scatter_req_0;
      aggregated_sig <= expr_645_wire_constant;
      array_obj_ref_644_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_648_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_648_gather_scatter_ack_0 <= array_obj_ref_648_gather_scatter_req_0;
      aggregated_sig <= expr_649_wire_constant;
      array_obj_ref_648_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_652_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_652_gather_scatter_ack_0 <= array_obj_ref_652_gather_scatter_req_0;
      aggregated_sig <= expr_653_wire_constant;
      array_obj_ref_652_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_656_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_656_gather_scatter_ack_0 <= array_obj_ref_656_gather_scatter_req_0;
      aggregated_sig <= expr_657_wire_constant;
      array_obj_ref_656_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_660_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_660_gather_scatter_ack_0 <= array_obj_ref_660_gather_scatter_req_0;
      aggregated_sig <= expr_661_wire_constant;
      array_obj_ref_660_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_664_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_664_gather_scatter_ack_0 <= array_obj_ref_664_gather_scatter_req_0;
      aggregated_sig <= expr_665_wire_constant;
      array_obj_ref_664_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_668_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_668_gather_scatter_ack_0 <= array_obj_ref_668_gather_scatter_req_0;
      aggregated_sig <= expr_669_wire_constant;
      array_obj_ref_668_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- shared store operator group (0) : array_obj_ref_640_store_0 array_obj_ref_636_store_0 array_obj_ref_644_store_0 array_obj_ref_648_store_0 array_obj_ref_652_store_0 array_obj_ref_656_store_0 array_obj_ref_660_store_0 array_obj_ref_664_store_0 array_obj_ref_668_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(35 downto 0);
      signal data_in: std_logic_vector(71 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 8 downto 0);
      -- 
    begin -- 
      reqL(8) <= array_obj_ref_640_store_0_req_0;
      reqL(7) <= array_obj_ref_636_store_0_req_0;
      reqL(6) <= array_obj_ref_644_store_0_req_0;
      reqL(5) <= array_obj_ref_648_store_0_req_0;
      reqL(4) <= array_obj_ref_652_store_0_req_0;
      reqL(3) <= array_obj_ref_656_store_0_req_0;
      reqL(2) <= array_obj_ref_660_store_0_req_0;
      reqL(1) <= array_obj_ref_664_store_0_req_0;
      reqL(0) <= array_obj_ref_668_store_0_req_0;
      array_obj_ref_640_store_0_ack_0 <= ackL(8);
      array_obj_ref_636_store_0_ack_0 <= ackL(7);
      array_obj_ref_644_store_0_ack_0 <= ackL(6);
      array_obj_ref_648_store_0_ack_0 <= ackL(5);
      array_obj_ref_652_store_0_ack_0 <= ackL(4);
      array_obj_ref_656_store_0_ack_0 <= ackL(3);
      array_obj_ref_660_store_0_ack_0 <= ackL(2);
      array_obj_ref_664_store_0_ack_0 <= ackL(1);
      array_obj_ref_668_store_0_ack_0 <= ackL(0);
      reqR(8) <= array_obj_ref_640_store_0_req_1;
      reqR(7) <= array_obj_ref_636_store_0_req_1;
      reqR(6) <= array_obj_ref_644_store_0_req_1;
      reqR(5) <= array_obj_ref_648_store_0_req_1;
      reqR(4) <= array_obj_ref_652_store_0_req_1;
      reqR(3) <= array_obj_ref_656_store_0_req_1;
      reqR(2) <= array_obj_ref_660_store_0_req_1;
      reqR(1) <= array_obj_ref_664_store_0_req_1;
      reqR(0) <= array_obj_ref_668_store_0_req_1;
      array_obj_ref_640_store_0_ack_1 <= ackR(8);
      array_obj_ref_636_store_0_ack_1 <= ackR(7);
      array_obj_ref_644_store_0_ack_1 <= ackR(6);
      array_obj_ref_648_store_0_ack_1 <= ackR(5);
      array_obj_ref_652_store_0_ack_1 <= ackR(4);
      array_obj_ref_656_store_0_ack_1 <= ackR(3);
      array_obj_ref_660_store_0_ack_1 <= ackR(2);
      array_obj_ref_664_store_0_ack_1 <= ackR(1);
      array_obj_ref_668_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_640_word_address_0 & array_obj_ref_636_word_address_0 & array_obj_ref_644_word_address_0 & array_obj_ref_648_word_address_0 & array_obj_ref_652_word_address_0 & array_obj_ref_656_word_address_0 & array_obj_ref_660_word_address_0 & array_obj_ref_664_word_address_0 & array_obj_ref_668_word_address_0;
      data_in <= array_obj_ref_640_data_0 & array_obj_ref_636_data_0 & array_obj_ref_644_data_0 & array_obj_ref_648_data_0 & array_obj_ref_652_data_0 & array_obj_ref_656_data_0 & array_obj_ref_660_data_0 & array_obj_ref_664_data_0 & array_obj_ref_668_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 9,
        tag_length => 4,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_11_sr_req(0),
          mack => memory_space_11_sr_ack(0),
          maddr => memory_space_11_sr_addr(3 downto 0),
          mdata => memory_space_11_sr_data(7 downto 0),
          mtag => memory_space_11_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 9,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_11_sc_req(0),
          mack => memory_space_11_sc_ack(0),
          mtag => memory_space_11_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity free_queue_manager is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(3 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(3 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(3 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(3 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(7 downto 0);
    free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_ack_pipe_write_data : out  std_logic_vector(7 downto 0);
    free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
    global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity free_queue_manager;
architecture Default of free_queue_manager is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal free_queue_manager_CP_3084_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_772_addr_0_ack_0 : boolean;
  signal ptr_deref_772_addr_0_req_0 : boolean;
  signal switch_stmt_730_branch_1_ack_1 : boolean;
  signal array_obj_ref_767_index_0_rename_req_0 : boolean;
  signal call_stmt_674_call_req_0 : boolean;
  signal binary_778_inst_req_1 : boolean;
  signal ptr_deref_693_gather_scatter_ack_0 : boolean;
  signal ptr_deref_682_store_0_req_1 : boolean;
  signal addr_of_768_final_reg_ack_0 : boolean;
  signal binary_778_inst_req_0 : boolean;
  signal binary_756_inst_ack_0 : boolean;
  signal ptr_deref_772_load_0_ack_1 : boolean;
  signal ptr_deref_693_store_0_req_0 : boolean;
  signal ptr_deref_772_base_resize_req_0 : boolean;
  signal call_stmt_674_call_ack_0 : boolean;
  signal switch_stmt_730_select_expr_0_req_0 : boolean;
  signal simple_obj_ref_728_inst_ack_0 : boolean;
  signal ptr_deref_693_gather_scatter_req_0 : boolean;
  signal switch_stmt_730_select_expr_1_ack_1 : boolean;
  signal switch_stmt_730_select_expr_1_req_1 : boolean;
  signal ptr_deref_704_gather_scatter_ack_0 : boolean;
  signal binary_791_inst_ack_0 : boolean;
  signal ptr_deref_772_load_0_req_1 : boolean;
  signal ptr_deref_772_base_resize_ack_0 : boolean;
  signal simple_obj_ref_728_inst_req_0 : boolean;
  signal binary_778_inst_ack_0 : boolean;
  signal switch_stmt_730_select_expr_0_ack_0 : boolean;
  signal ptr_deref_682_store_0_ack_1 : boolean;
  signal array_obj_ref_767_offset_inst_req_0 : boolean;
  signal if_stmt_758_branch_ack_0 : boolean;
  signal switch_stmt_730_select_expr_1_req_0 : boolean;
  signal binary_756_inst_req_0 : boolean;
  signal switch_stmt_730_branch_default_ack_0 : boolean;
  signal switch_stmt_730_branch_1_req_0 : boolean;
  signal binary_778_inst_ack_1 : boolean;
  signal type_cast_752_inst_ack_0 : boolean;
  signal ptr_deref_693_store_0_ack_0 : boolean;
  signal ptr_deref_715_store_0_req_0 : boolean;
  signal if_stmt_780_branch_req_0 : boolean;
  signal ptr_deref_772_gather_scatter_req_0 : boolean;
  signal binary_756_inst_ack_1 : boolean;
  signal ptr_deref_704_store_0_ack_1 : boolean;
  signal addr_of_768_final_reg_req_0 : boolean;
  signal binary_756_inst_req_1 : boolean;
  signal switch_stmt_730_branch_0_ack_1 : boolean;
  signal binary_791_inst_req_0 : boolean;
  signal ptr_deref_682_gather_scatter_ack_0 : boolean;
  signal if_stmt_758_branch_req_0 : boolean;
  signal switch_stmt_730_select_expr_1_ack_0 : boolean;
  signal ptr_deref_715_store_0_ack_1 : boolean;
  signal ptr_deref_693_store_0_req_1 : boolean;
  signal type_cast_752_inst_req_0 : boolean;
  signal array_obj_ref_767_index_0_resize_req_0 : boolean;
  signal array_obj_ref_767_index_0_rename_ack_0 : boolean;
  signal switch_stmt_730_branch_0_req_0 : boolean;
  signal ptr_deref_715_store_0_req_1 : boolean;
  signal ptr_deref_704_gather_scatter_req_0 : boolean;
  signal ptr_deref_682_store_0_ack_0 : boolean;
  signal ptr_deref_715_store_0_ack_0 : boolean;
  signal ptr_deref_693_store_0_ack_1 : boolean;
  signal ptr_deref_704_store_0_req_0 : boolean;
  signal switch_stmt_730_select_expr_0_req_1 : boolean;
  signal if_stmt_758_branch_ack_1 : boolean;
  signal ptr_deref_682_store_0_req_0 : boolean;
  signal ptr_deref_715_gather_scatter_ack_0 : boolean;
  signal ptr_deref_772_load_0_ack_0 : boolean;
  signal ptr_deref_715_gather_scatter_req_0 : boolean;
  signal switch_stmt_730_select_expr_0_ack_1 : boolean;
  signal ptr_deref_772_root_address_inst_req_0 : boolean;
  signal array_obj_ref_767_root_address_inst_req_0 : boolean;
  signal ptr_deref_772_load_0_req_0 : boolean;
  signal array_obj_ref_767_offset_inst_ack_0 : boolean;
  signal if_stmt_780_branch_ack_0 : boolean;
  signal ptr_deref_704_store_0_req_1 : boolean;
  signal binary_791_inst_ack_1 : boolean;
  signal switch_stmt_730_branch_default_req_0 : boolean;
  signal ptr_deref_682_gather_scatter_req_0 : boolean;
  signal binary_791_inst_req_1 : boolean;
  signal array_obj_ref_767_index_0_resize_ack_0 : boolean;
  signal call_stmt_674_call_req_1 : boolean;
  signal call_stmt_674_call_ack_1 : boolean;
  signal ptr_deref_772_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_767_root_address_inst_ack_0 : boolean;
  signal ptr_deref_772_gather_scatter_ack_0 : boolean;
  signal if_stmt_780_branch_ack_1 : boolean;
  signal array_obj_ref_803_root_address_inst_req_0 : boolean;
  signal array_obj_ref_803_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_803_root_address_inst_req_1 : boolean;
  signal array_obj_ref_803_root_address_inst_ack_1 : boolean;
  signal ptr_deref_811_base_resize_req_0 : boolean;
  signal ptr_deref_811_base_resize_ack_0 : boolean;
  signal array_obj_ref_803_offset_inst_ack_0 : boolean;
  signal array_obj_ref_803_offset_inst_req_0 : boolean;
  signal array_obj_ref_803_index_0_rename_req_0 : boolean;
  signal array_obj_ref_803_index_0_rename_ack_0 : boolean;
  signal type_cast_808_inst_req_0 : boolean;
  signal type_cast_808_inst_ack_0 : boolean;
  signal array_obj_ref_803_index_0_resize_req_0 : boolean;
  signal array_obj_ref_803_index_0_resize_ack_0 : boolean;
  signal addr_of_804_final_reg_ack_0 : boolean;
  signal binary_799_inst_ack_1 : boolean;
  signal addr_of_804_final_reg_req_0 : boolean;
  signal binary_799_inst_ack_0 : boolean;
  signal binary_799_inst_req_1 : boolean;
  signal ptr_deref_811_root_address_inst_req_0 : boolean;
  signal ptr_deref_811_root_address_inst_ack_0 : boolean;
  signal binary_799_inst_req_0 : boolean;
  signal ptr_deref_704_store_0_ack_0 : boolean;
  signal ptr_deref_811_addr_0_req_0 : boolean;
  signal ptr_deref_811_addr_0_ack_0 : boolean;
  signal ptr_deref_811_gather_scatter_req_0 : boolean;
  signal ptr_deref_811_gather_scatter_ack_0 : boolean;
  signal ptr_deref_811_store_0_req_0 : boolean;
  signal ptr_deref_811_store_0_ack_0 : boolean;
  signal ptr_deref_811_store_0_req_1 : boolean;
  signal ptr_deref_811_store_0_ack_1 : boolean;
  signal simple_obj_ref_821_inst_req_0 : boolean;
  signal simple_obj_ref_821_inst_ack_0 : boolean;
  signal simple_obj_ref_831_inst_req_0 : boolean;
  signal simple_obj_ref_831_inst_ack_0 : boolean;
  signal simple_obj_ref_842_inst_req_0 : boolean;
  signal simple_obj_ref_842_inst_ack_0 : boolean;
  signal simple_obj_ref_855_inst_req_0 : boolean;
  signal simple_obj_ref_855_inst_ack_0 : boolean;
  signal binary_861_inst_req_0 : boolean;
  signal binary_861_inst_ack_0 : boolean;
  signal binary_861_inst_req_1 : boolean;
  signal binary_861_inst_ack_1 : boolean;
  signal if_stmt_863_branch_req_0 : boolean;
  signal if_stmt_863_branch_ack_1 : boolean;
  signal if_stmt_863_branch_ack_0 : boolean;
  signal binary_882_inst_req_0 : boolean;
  signal binary_882_inst_ack_0 : boolean;
  signal binary_882_inst_req_1 : boolean;
  signal binary_882_inst_ack_1 : boolean;
  signal binary_888_inst_req_0 : boolean;
  signal binary_888_inst_ack_0 : boolean;
  signal binary_888_inst_req_1 : boolean;
  signal binary_888_inst_ack_1 : boolean;
  signal binary_894_inst_req_0 : boolean;
  signal binary_894_inst_ack_0 : boolean;
  signal binary_894_inst_req_1 : boolean;
  signal binary_894_inst_ack_1 : boolean;
  signal binary_899_inst_req_0 : boolean;
  signal binary_899_inst_ack_0 : boolean;
  signal binary_899_inst_req_1 : boolean;
  signal binary_899_inst_ack_1 : boolean;
  signal if_stmt_901_branch_req_0 : boolean;
  signal if_stmt_901_branch_ack_1 : boolean;
  signal if_stmt_901_branch_ack_0 : boolean;
  signal type_cast_910_inst_req_0 : boolean;
  signal type_cast_910_inst_ack_0 : boolean;
  signal binary_914_inst_req_0 : boolean;
  signal binary_914_inst_ack_0 : boolean;
  signal binary_914_inst_req_1 : boolean;
  signal binary_914_inst_ack_1 : boolean;
  signal if_stmt_916_branch_req_0 : boolean;
  signal if_stmt_916_branch_ack_1 : boolean;
  signal if_stmt_916_branch_ack_0 : boolean;
  signal array_obj_ref_933_index_0_resize_req_0 : boolean;
  signal array_obj_ref_933_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_933_index_0_rename_req_0 : boolean;
  signal array_obj_ref_933_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_933_offset_inst_req_0 : boolean;
  signal array_obj_ref_933_offset_inst_ack_0 : boolean;
  signal array_obj_ref_933_root_address_inst_req_0 : boolean;
  signal array_obj_ref_933_root_address_inst_ack_0 : boolean;
  signal addr_of_934_final_reg_req_0 : boolean;
  signal addr_of_934_final_reg_ack_0 : boolean;
  signal ptr_deref_937_base_resize_req_0 : boolean;
  signal ptr_deref_937_base_resize_ack_0 : boolean;
  signal ptr_deref_937_root_address_inst_req_0 : boolean;
  signal ptr_deref_937_root_address_inst_ack_0 : boolean;
  signal ptr_deref_937_addr_0_req_0 : boolean;
  signal ptr_deref_937_addr_0_ack_0 : boolean;
  signal ptr_deref_937_gather_scatter_req_0 : boolean;
  signal ptr_deref_937_gather_scatter_ack_0 : boolean;
  signal ptr_deref_937_store_0_req_0 : boolean;
  signal ptr_deref_937_store_0_ack_0 : boolean;
  signal ptr_deref_937_store_0_req_1 : boolean;
  signal ptr_deref_937_store_0_ack_1 : boolean;
  signal type_cast_744_inst_req_0 : boolean;
  signal type_cast_744_inst_ack_0 : boolean;
  signal phi_stmt_741_req_0 : boolean;
  signal phi_stmt_741_req_1 : boolean;
  signal phi_stmt_741_ack_0 : boolean;
  signal phi_stmt_870_req_1 : boolean;
  signal type_cast_873_inst_req_0 : boolean;
  signal type_cast_873_inst_ack_0 : boolean;
  signal phi_stmt_870_req_0 : boolean;
  signal phi_stmt_870_ack_0 : boolean;
  signal phi_stmt_923_req_1 : boolean;
  signal type_cast_926_inst_req_0 : boolean;
  signal type_cast_926_inst_ack_0 : boolean;
  signal phi_stmt_923_req_0 : boolean;
  signal phi_stmt_923_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  free_queue_manager_CP_3084: Block -- control-path 
    signal cp_elements: BooleanArray(258 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    call_stmt_674_call_req_0 <= cp_elements(0);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(45);
    cp_elements(3) <= OrReduce(cp_elements(236) & cp_elements(240));
    cp_elements(4) <= OrReduce(cp_elements(81) & cp_elements(242));
    cp_elements(5) <= OrReduce(cp_elements(113) & cp_elements(244));
    cp_elements(6) <= cp_elements(147);
    simple_obj_ref_821_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= OrReduce(cp_elements(246) & cp_elements(250));
    cp_elements(8) <= cp_elements(187);
    cp_elements(9) <= OrReduce(cp_elements(196) & cp_elements(252));
    cp_elements(10) <= OrReduce(cp_elements(254) & cp_elements(258));
    cp_elements(11) <= call_stmt_674_call_ack_0;
    call_stmt_674_call_req_1 <= cp_elements(11);
    cp_elements(12) <= call_stmt_674_call_ack_1;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= cp_elements(13);
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(17));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_682_gather_scatter_req_0 <= cp_elements(15);
    cp_elements(16) <= cp_elements(13);
    cp_elements(17) <= cp_elements(13);
    cp_elements(18) <= ptr_deref_682_gather_scatter_ack_0;
    ptr_deref_682_store_0_req_0 <= cp_elements(18);
    cp_elements(19) <= ptr_deref_682_store_0_ack_0;
    cp_elements(20) <= cp_elements(19);
    ptr_deref_682_store_0_req_1 <= cp_elements(20);
    cp_elements(21) <= ptr_deref_682_store_0_ack_1;
    cp_elements(22) <= cp_elements(13);
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(22) & cp_elements(25));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_693_gather_scatter_req_0 <= cp_elements(23);
    cp_elements(24) <= cp_elements(13);
    cp_elements(25) <= cp_elements(13);
    cp_elements(26) <= ptr_deref_693_gather_scatter_ack_0;
    ptr_deref_693_store_0_req_0 <= cp_elements(26);
    cp_elements(27) <= ptr_deref_693_store_0_ack_0;
    cp_elements(28) <= cp_elements(27);
    ptr_deref_693_store_0_req_1 <= cp_elements(28);
    cp_elements(29) <= ptr_deref_693_store_0_ack_1;
    cp_elements(30) <= cp_elements(13);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(30) & cp_elements(33));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_704_gather_scatter_req_0 <= cp_elements(31);
    cp_elements(32) <= cp_elements(13);
    cp_elements(33) <= cp_elements(13);
    cp_elements(34) <= ptr_deref_704_gather_scatter_ack_0;
    ptr_deref_704_store_0_req_0 <= cp_elements(34);
    cp_elements(35) <= ptr_deref_704_store_0_ack_0;
    cp_elements(36) <= cp_elements(35);
    ptr_deref_704_store_0_req_1 <= cp_elements(36);
    cp_elements(37) <= ptr_deref_704_store_0_ack_1;
    cp_elements(38) <= cp_elements(13);
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38) & cp_elements(41));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_715_gather_scatter_req_0 <= cp_elements(39);
    cp_elements(40) <= cp_elements(13);
    cp_elements(41) <= cp_elements(13);
    cp_elements(42) <= ptr_deref_715_gather_scatter_ack_0;
    ptr_deref_715_store_0_req_0 <= cp_elements(42);
    cp_elements(43) <= ptr_deref_715_store_0_ack_0;
    ptr_deref_715_store_0_req_1 <= cp_elements(43);
    cp_elements(44) <= ptr_deref_715_store_0_ack_1;
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(21) & cp_elements(24) & cp_elements(29) & cp_elements(32) & cp_elements(37) & cp_elements(40) & cp_elements(44));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= simple_obj_ref_728_inst_ack_0;
    cp_elements(47) <= cp_elements(46);
    cp_elements(48) <= false;
    cp_elements(49) <= cp_elements(48);
    cp_elements(50) <= cp_elements(46);
    cp_elements(51) <= cp_elements(50);
    cp_elements(52) <= cp_elements(51);
    switch_stmt_730_select_expr_0_req_0 <= cp_elements(52);
    cp_elements(53) <= switch_stmt_730_select_expr_0_ack_0;
    switch_stmt_730_select_expr_0_req_1 <= cp_elements(53);
    cp_elements(54) <= switch_stmt_730_select_expr_0_ack_1;
    switch_stmt_730_branch_0_req_0 <= cp_elements(54);
    cp_elements(55) <= cp_elements(51);
    switch_stmt_730_select_expr_1_req_0 <= cp_elements(55);
    cp_elements(56) <= switch_stmt_730_select_expr_1_ack_0;
    switch_stmt_730_select_expr_1_req_1 <= cp_elements(56);
    cp_elements(57) <= switch_stmt_730_select_expr_1_ack_1;
    switch_stmt_730_branch_1_req_0 <= cp_elements(57);
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(54) & cp_elements(57));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    switch_stmt_730_branch_default_req_0 <= cp_elements(58);
    cp_elements(59) <= cp_elements(58);
    cp_elements(60) <= cp_elements(59);
    cp_elements(61) <= switch_stmt_730_branch_0_ack_1;
    phi_stmt_741_req_1 <= cp_elements(61);
    cp_elements(62) <= cp_elements(59);
    cp_elements(63) <= switch_stmt_730_branch_1_ack_1;
    simple_obj_ref_855_inst_req_0 <= cp_elements(63);
    cp_elements(64) <= cp_elements(59);
    cp_elements(65) <= switch_stmt_730_branch_default_ack_0;
    cp_elements(66) <= cp_elements(3);
    cpelement_group_67 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(72));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(67),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_756_inst_req_0 <= cp_elements(67);
    cp_elements(68) <= cp_elements(66);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(70) & cp_elements(71));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_752_inst_req_0 <= cp_elements(69);
    cp_elements(70) <= cp_elements(66);
    cp_elements(71) <= cp_elements(66);
    cp_elements(72) <= type_cast_752_inst_ack_0;
    cp_elements(73) <= binary_756_inst_ack_0;
    binary_756_inst_req_1 <= cp_elements(73);
    cp_elements(74) <= binary_756_inst_ack_1;
    cp_elements(75) <= cp_elements(74);
    cp_elements(76) <= false;
    cp_elements(77) <= cp_elements(76);
    cp_elements(78) <= cp_elements(74);
    if_stmt_758_branch_req_0 <= cp_elements(78);
    cp_elements(79) <= cp_elements(78);
    cp_elements(80) <= cp_elements(79);
    cp_elements(81) <= if_stmt_758_branch_ack_1;
    cp_elements(82) <= cp_elements(79);
    cp_elements(83) <= if_stmt_758_branch_ack_0;
    simple_obj_ref_842_inst_req_0 <= cp_elements(83);
    cp_elements(84) <= cp_elements(4);
    cpelement_group_85 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(86) & cp_elements(91));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(85),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_768_final_reg_req_0 <= cp_elements(85);
    cp_elements(86) <= cp_elements(84);
    cp_elements(87) <= cp_elements(84);
    array_obj_ref_767_index_0_resize_req_0 <= cp_elements(87);
    cp_elements(88) <= array_obj_ref_767_index_0_resize_ack_0;
    array_obj_ref_767_index_0_rename_req_0 <= cp_elements(88);
    cp_elements(89) <= array_obj_ref_767_index_0_rename_ack_0;
    array_obj_ref_767_offset_inst_req_0 <= cp_elements(89);
    cp_elements(90) <= array_obj_ref_767_offset_inst_ack_0;
    array_obj_ref_767_root_address_inst_req_0 <= cp_elements(90);
    cp_elements(91) <= array_obj_ref_767_root_address_inst_ack_0;
    cp_elements(92) <= addr_of_768_final_reg_ack_0;
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(92) & cp_elements(97));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_772_load_0_req_0 <= cp_elements(93);
    cp_elements(94) <= cp_elements(92);
    ptr_deref_772_base_resize_req_0 <= cp_elements(94);
    cp_elements(95) <= ptr_deref_772_base_resize_ack_0;
    ptr_deref_772_root_address_inst_req_0 <= cp_elements(95);
    cp_elements(96) <= ptr_deref_772_root_address_inst_ack_0;
    ptr_deref_772_addr_0_req_0 <= cp_elements(96);
    cp_elements(97) <= ptr_deref_772_addr_0_ack_0;
    cp_elements(98) <= ptr_deref_772_load_0_ack_0;
    ptr_deref_772_load_0_req_1 <= cp_elements(98);
    cp_elements(99) <= ptr_deref_772_load_0_ack_1;
    ptr_deref_772_gather_scatter_req_0 <= cp_elements(99);
    cp_elements(100) <= ptr_deref_772_gather_scatter_ack_0;
    cpelement_group_101 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(100) & cp_elements(102));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(101),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_778_inst_req_0 <= cp_elements(101);
    cp_elements(102) <= cp_elements(84);
    cp_elements(103) <= binary_778_inst_ack_0;
    binary_778_inst_req_1 <= cp_elements(103);
    cp_elements(104) <= binary_778_inst_ack_1;
    cp_elements(105) <= cp_elements(104);
    cp_elements(106) <= false;
    cp_elements(107) <= cp_elements(106);
    cp_elements(108) <= cp_elements(104);
    if_stmt_780_branch_req_0 <= cp_elements(108);
    cp_elements(109) <= cp_elements(108);
    cp_elements(110) <= cp_elements(109);
    cp_elements(111) <= if_stmt_780_branch_ack_1;
    cp_elements(112) <= cp_elements(109);
    cp_elements(113) <= if_stmt_780_branch_ack_0;
    cp_elements(114) <= cp_elements(5);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(116) & cp_elements(117));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_791_inst_req_0 <= cp_elements(115);
    cp_elements(116) <= cp_elements(114);
    cp_elements(117) <= cp_elements(114);
    cp_elements(118) <= binary_791_inst_ack_0;
    binary_791_inst_req_1 <= cp_elements(118);
    cp_elements(119) <= binary_791_inst_ack_1;
    type_cast_744_inst_req_0 <= cp_elements(119);
    cp_elements(120) <= cp_elements(111);
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(122) & cp_elements(123));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_799_inst_req_0 <= cp_elements(121);
    cp_elements(122) <= cp_elements(120);
    cp_elements(123) <= cp_elements(120);
    cp_elements(124) <= binary_799_inst_ack_0;
    binary_799_inst_req_1 <= cp_elements(124);
    cp_elements(125) <= binary_799_inst_ack_1;
    array_obj_ref_803_index_0_resize_req_0 <= cp_elements(125);
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(132));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_804_final_reg_req_0 <= cp_elements(126);
    cp_elements(127) <= cp_elements(120);
    cp_elements(128) <= array_obj_ref_803_index_0_resize_ack_0;
    array_obj_ref_803_index_0_rename_req_0 <= cp_elements(128);
    cp_elements(129) <= array_obj_ref_803_index_0_rename_ack_0;
    array_obj_ref_803_offset_inst_req_0 <= cp_elements(129);
    cp_elements(130) <= array_obj_ref_803_offset_inst_ack_0;
    array_obj_ref_803_root_address_inst_req_0 <= cp_elements(130);
    cp_elements(131) <= array_obj_ref_803_root_address_inst_ack_0;
    array_obj_ref_803_root_address_inst_req_1 <= cp_elements(131);
    cp_elements(132) <= array_obj_ref_803_root_address_inst_ack_1;
    cp_elements(133) <= addr_of_804_final_reg_ack_0;
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(133) & cp_elements(135));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_808_inst_req_0 <= cp_elements(134);
    cp_elements(135) <= cp_elements(120);
    cp_elements(136) <= type_cast_808_inst_ack_0;
    cp_elements(137) <= cp_elements(120);
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(139) & cp_elements(143));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_811_gather_scatter_req_0 <= cp_elements(138);
    cp_elements(139) <= cp_elements(120);
    cp_elements(140) <= cp_elements(139);
    ptr_deref_811_base_resize_req_0 <= cp_elements(140);
    cp_elements(141) <= ptr_deref_811_base_resize_ack_0;
    ptr_deref_811_root_address_inst_req_0 <= cp_elements(141);
    cp_elements(142) <= ptr_deref_811_root_address_inst_ack_0;
    ptr_deref_811_addr_0_req_0 <= cp_elements(142);
    cp_elements(143) <= ptr_deref_811_addr_0_ack_0;
    cp_elements(144) <= ptr_deref_811_gather_scatter_ack_0;
    ptr_deref_811_store_0_req_0 <= cp_elements(144);
    cp_elements(145) <= ptr_deref_811_store_0_ack_0;
    ptr_deref_811_store_0_req_1 <= cp_elements(145);
    cp_elements(146) <= ptr_deref_811_store_0_ack_1;
    cpelement_group_147 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(136) & cp_elements(146));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(148) <= simple_obj_ref_821_inst_ack_0;
    simple_obj_ref_831_inst_req_0 <= cp_elements(148);
    cp_elements(149) <= simple_obj_ref_831_inst_ack_0;
    cp_elements(150) <= simple_obj_ref_842_inst_ack_0;
    cp_elements(151) <= simple_obj_ref_855_inst_ack_0;
    cp_elements(152) <= cp_elements(151);
    cpelement_group_153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(154) & cp_elements(155));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_861_inst_req_0 <= cp_elements(153);
    cp_elements(154) <= cp_elements(152);
    cp_elements(155) <= cp_elements(152);
    cp_elements(156) <= binary_861_inst_ack_0;
    binary_861_inst_req_1 <= cp_elements(156);
    cp_elements(157) <= binary_861_inst_ack_1;
    cp_elements(158) <= cp_elements(157);
    cp_elements(159) <= false;
    cp_elements(160) <= cp_elements(159);
    cp_elements(161) <= cp_elements(157);
    if_stmt_863_branch_req_0 <= cp_elements(161);
    cp_elements(162) <= cp_elements(161);
    cp_elements(163) <= cp_elements(162);
    cp_elements(164) <= if_stmt_863_branch_ack_1;
    phi_stmt_870_req_1 <= cp_elements(164);
    cp_elements(165) <= cp_elements(162);
    cp_elements(166) <= if_stmt_863_branch_ack_0;
    phi_stmt_923_req_1 <= cp_elements(166);
    cp_elements(167) <= cp_elements(7);
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_882_inst_req_0 <= cp_elements(168);
    cp_elements(169) <= cp_elements(167);
    cp_elements(170) <= cp_elements(167);
    cp_elements(171) <= binary_882_inst_ack_0;
    binary_882_inst_req_1 <= cp_elements(171);
    cp_elements(172) <= binary_882_inst_ack_1;
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(174) & cp_elements(175));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_888_inst_req_0 <= cp_elements(173);
    cp_elements(174) <= cp_elements(167);
    cp_elements(175) <= cp_elements(167);
    cp_elements(176) <= binary_888_inst_ack_0;
    binary_888_inst_req_1 <= cp_elements(176);
    cp_elements(177) <= binary_888_inst_ack_1;
    cpelement_group_178 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(179));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(178),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_894_inst_req_0 <= cp_elements(178);
    cp_elements(179) <= cp_elements(167);
    cp_elements(180) <= binary_894_inst_ack_0;
    binary_894_inst_req_1 <= cp_elements(180);
    cp_elements(181) <= binary_894_inst_ack_1;
    cpelement_group_182 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(183) & cp_elements(184));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(182),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_899_inst_req_0 <= cp_elements(182);
    cp_elements(183) <= cp_elements(167);
    cp_elements(184) <= cp_elements(167);
    cp_elements(185) <= binary_899_inst_ack_0;
    binary_899_inst_req_1 <= cp_elements(185);
    cp_elements(186) <= binary_899_inst_ack_1;
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(177) & cp_elements(186));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(188) <= cp_elements(8);
    cp_elements(189) <= false;
    cp_elements(190) <= cp_elements(189);
    cp_elements(191) <= cp_elements(8);
    if_stmt_901_branch_req_0 <= cp_elements(191);
    cp_elements(192) <= cp_elements(191);
    cp_elements(193) <= cp_elements(192);
    cp_elements(194) <= if_stmt_901_branch_ack_1;
    type_cast_873_inst_req_0 <= cp_elements(194);
    cp_elements(195) <= cp_elements(192);
    cp_elements(196) <= if_stmt_901_branch_ack_0;
    cp_elements(197) <= cp_elements(9);
    cpelement_group_198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(199) & cp_elements(203));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_914_inst_req_0 <= cp_elements(198);
    cp_elements(199) <= cp_elements(197);
    cpelement_group_200 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(201) & cp_elements(202));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(200),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_910_inst_req_0 <= cp_elements(200);
    cp_elements(201) <= cp_elements(197);
    cp_elements(202) <= cp_elements(197);
    cp_elements(203) <= type_cast_910_inst_ack_0;
    cp_elements(204) <= binary_914_inst_ack_0;
    binary_914_inst_req_1 <= cp_elements(204);
    cp_elements(205) <= binary_914_inst_ack_1;
    cp_elements(206) <= cp_elements(205);
    cp_elements(207) <= false;
    cp_elements(208) <= cp_elements(207);
    cp_elements(209) <= cp_elements(205);
    if_stmt_916_branch_req_0 <= cp_elements(209);
    cp_elements(210) <= cp_elements(209);
    cp_elements(211) <= cp_elements(210);
    cp_elements(212) <= if_stmt_916_branch_ack_1;
    type_cast_926_inst_req_0 <= cp_elements(212);
    cp_elements(213) <= cp_elements(210);
    cp_elements(214) <= if_stmt_916_branch_ack_0;
    cp_elements(215) <= cp_elements(10);
    cpelement_group_216 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(217) & cp_elements(222));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(216),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_934_final_reg_req_0 <= cp_elements(216);
    cp_elements(217) <= cp_elements(215);
    cp_elements(218) <= cp_elements(215);
    array_obj_ref_933_index_0_resize_req_0 <= cp_elements(218);
    cp_elements(219) <= array_obj_ref_933_index_0_resize_ack_0;
    array_obj_ref_933_index_0_rename_req_0 <= cp_elements(219);
    cp_elements(220) <= array_obj_ref_933_index_0_rename_ack_0;
    array_obj_ref_933_offset_inst_req_0 <= cp_elements(220);
    cp_elements(221) <= array_obj_ref_933_offset_inst_ack_0;
    array_obj_ref_933_root_address_inst_req_0 <= cp_elements(221);
    cp_elements(222) <= array_obj_ref_933_root_address_inst_ack_0;
    cp_elements(223) <= addr_of_934_final_reg_ack_0;
    cp_elements(224) <= cp_elements(215);
    cpelement_group_225 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(224) & cp_elements(229));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(225),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_937_gather_scatter_req_0 <= cp_elements(225);
    cp_elements(226) <= cp_elements(223);
    ptr_deref_937_base_resize_req_0 <= cp_elements(226);
    cp_elements(227) <= ptr_deref_937_base_resize_ack_0;
    ptr_deref_937_root_address_inst_req_0 <= cp_elements(227);
    cp_elements(228) <= ptr_deref_937_root_address_inst_ack_0;
    ptr_deref_937_addr_0_req_0 <= cp_elements(228);
    cp_elements(229) <= ptr_deref_937_addr_0_ack_0;
    cp_elements(230) <= ptr_deref_937_gather_scatter_ack_0;
    ptr_deref_937_store_0_req_0 <= cp_elements(230);
    cp_elements(231) <= ptr_deref_937_store_0_ack_0;
    ptr_deref_937_store_0_req_1 <= cp_elements(231);
    cp_elements(232) <= ptr_deref_937_store_0_ack_1;
    cp_elements(233) <= OrReduce(cp_elements(2) & cp_elements(65) & cp_elements(149) & cp_elements(150) & cp_elements(214) & cp_elements(232));
    cp_elements(234) <= cp_elements(233);
    simple_obj_ref_728_inst_req_0 <= cp_elements(234);
    cp_elements(235) <= false;
    cp_elements(236) <= cp_elements(235);
    cp_elements(237) <= type_cast_744_inst_ack_0;
    phi_stmt_741_req_0 <= cp_elements(237);
    cp_elements(238) <= OrReduce(cp_elements(61) & cp_elements(237));
    cp_elements(239) <= cp_elements(238);
    cp_elements(240) <= phi_stmt_741_ack_0;
    cp_elements(241) <= false;
    cp_elements(242) <= cp_elements(241);
    cp_elements(243) <= false;
    cp_elements(244) <= cp_elements(243);
    cp_elements(245) <= false;
    cp_elements(246) <= cp_elements(245);
    cp_elements(247) <= type_cast_873_inst_ack_0;
    phi_stmt_870_req_0 <= cp_elements(247);
    cp_elements(248) <= OrReduce(cp_elements(164) & cp_elements(247));
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= phi_stmt_870_ack_0;
    cp_elements(251) <= false;
    cp_elements(252) <= cp_elements(251);
    cp_elements(253) <= false;
    cp_elements(254) <= cp_elements(253);
    cp_elements(255) <= type_cast_926_inst_ack_0;
    phi_stmt_923_req_0 <= cp_elements(255);
    cp_elements(256) <= OrReduce(cp_elements(166) & cp_elements(255));
    cp_elements(257) <= cp_elements(256);
    cp_elements(258) <= phi_stmt_923_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_767_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_767_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_767_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_767_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_803_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_803_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_803_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_803_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_933_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_933_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_933_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_933_root_address : std_logic_vector(2 downto 0);
    signal expr_732_wire_constant : std_logic_vector(7 downto 0);
    signal expr_732_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_735_wire_constant : std_logic_vector(7 downto 0);
    signal expr_735_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal i3x_x044_870 : std_logic_vector(31 downto 0);
    signal i3x_x0x_xlcssa53_923 : std_logic_vector(31 downto 0);
    signal iNsTr_10_726 : std_logic_vector(31 downto 0);
    signal iNsTr_12_741 : std_logic_vector(31 downto 0);
    signal iNsTr_14_853 : std_logic_vector(31 downto 0);
    signal iNsTr_17_841 : std_logic_vector(31 downto 0);
    signal iNsTr_1_680 : std_logic_vector(31 downto 0);
    signal iNsTr_20_889 : std_logic_vector(31 downto 0);
    signal iNsTr_25_820 : std_logic_vector(31 downto 0);
    signal iNsTr_27_830 : std_logic_vector(31 downto 0);
    signal iNsTr_3_691 : std_logic_vector(31 downto 0);
    signal iNsTr_5_702 : std_logic_vector(31 downto 0);
    signal iNsTr_7_713 : std_logic_vector(31 downto 0);
    signal ptr_deref_682_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_682_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_682_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_693_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_693_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_693_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_704_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_704_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_704_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_715_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_715_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_715_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_772_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_772_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_772_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_772_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_772_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_811_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_811_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_811_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_811_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_811_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_811_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_937_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_937_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_937_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_937_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_937_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_937_word_offset_0 : std_logic_vector(2 downto 0);
    signal simple_obj_ref_766_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_766_scaled : std_logic_vector(2 downto 0);
    signal simple_obj_ref_802_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_802_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_932_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_932_scaled : std_logic_vector(2 downto 0);
    signal tmp10_757 : std_logic_vector(0 downto 0);
    signal tmp12_769 : std_logic_vector(31 downto 0);
    signal tmp13_773 : std_logic_vector(7 downto 0);
    signal tmp14_779 : std_logic_vector(0 downto 0);
    signal tmp16_800 : std_logic_vector(31 downto 0);
    signal tmp17_805 : std_logic_vector(31 downto 0);
    signal tmp18_809 : std_logic_vector(31 downto 0);
    signal tmp21_792 : std_logic_vector(31 downto 0);
    signal tmp28_856 : std_logic_vector(31 downto 0);
    signal tmp31_895 : std_logic_vector(31 downto 0);
    signal tmp3243_862 : std_logic_vector(0 downto 0);
    signal tmp32_900 : std_logic_vector(0 downto 0);
    signal tmp36_915 : std_logic_vector(0 downto 0);
    signal tmp38_935 : std_logic_vector(31 downto 0);
    signal tmp50_883 : std_logic_vector(31 downto 0);
    signal tmp6_729 : std_logic_vector(7 downto 0);
    signal type_cast_684_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_695_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_706_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_717_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_744_wire : std_logic_vector(31 downto 0);
    signal type_cast_747_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_752_wire : std_logic_vector(31 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_777_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_790_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_798_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_813_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_823_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_844_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_860_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_873_wire : std_logic_vector(31 downto 0);
    signal type_cast_876_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_881_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_887_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_910_wire : std_logic_vector(31 downto 0);
    signal type_cast_913_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_926_wire : std_logic_vector(31 downto 0);
    signal type_cast_929_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_939_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_767_offset_scale_factor_0 <= "001";
    array_obj_ref_767_resized_base_address <= "000";
    array_obj_ref_803_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_803_resized_base_address <= "00000000001";
    array_obj_ref_933_offset_scale_factor_0 <= "001";
    array_obj_ref_933_resized_base_address <= "000";
    expr_732_wire_constant <= "00000010";
    expr_735_wire_constant <= "00000001";
    iNsTr_10_726 <= "00000000000000000000000000000000";
    iNsTr_14_853 <= "00000000000000000000000000000000";
    iNsTr_17_841 <= "00000000000000000000000000000000";
    iNsTr_1_680 <= "00000000000000000000000000000000";
    iNsTr_25_820 <= "00000000000000000000000000000000";
    iNsTr_27_830 <= "00000000000000000000000000000000";
    iNsTr_3_691 <= "00000000000000000000000000000001";
    iNsTr_5_702 <= "00000000000000000000000000000010";
    iNsTr_7_713 <= "00000000000000000000000000000011";
    ptr_deref_682_word_address_0 <= "000";
    ptr_deref_693_word_address_0 <= "001";
    ptr_deref_704_word_address_0 <= "010";
    ptr_deref_715_word_address_0 <= "011";
    ptr_deref_772_word_offset_0 <= "000";
    ptr_deref_811_word_offset_0 <= "000";
    ptr_deref_937_word_offset_0 <= "000";
    type_cast_684_wire_constant <= "00000001";
    type_cast_695_wire_constant <= "00000001";
    type_cast_706_wire_constant <= "00000001";
    type_cast_717_wire_constant <= "00000001";
    type_cast_747_wire_constant <= "00000000000000000000000000000000";
    type_cast_755_wire_constant <= "00000000000000000000000000000100";
    type_cast_777_wire_constant <= "00000001";
    type_cast_790_wire_constant <= "00000000000000000000000000000001";
    type_cast_798_wire_constant <= "00000000000000000000000000001000";
    type_cast_813_wire_constant <= "00000000";
    type_cast_823_wire_constant <= "00000011";
    type_cast_844_wire_constant <= "00000100";
    type_cast_860_wire_constant <= "00000000000000000000000100000000";
    type_cast_876_wire_constant <= "00000000000000000000000000000000";
    type_cast_881_wire_constant <= "00000000000000000000000000001000";
    type_cast_887_wire_constant <= "00000000000000000000000000000001";
    type_cast_893_wire_constant <= "00000000000000000000001000000000";
    type_cast_913_wire_constant <= "00000000000000000000000000000100";
    type_cast_929_wire_constant <= "00000000000000000000000000000000";
    type_cast_939_wire_constant <= "00000001";
    phi_stmt_741: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_744_wire & type_cast_747_wire_constant;
      req <= phi_stmt_741_req_0 & phi_stmt_741_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_741_ack_0,
          idata => idata,
          odata => iNsTr_12_741,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_741
    phi_stmt_870: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_873_wire & type_cast_876_wire_constant;
      req <= phi_stmt_870_req_0 & phi_stmt_870_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_870_ack_0,
          idata => idata,
          odata => i3x_x044_870,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_870
    phi_stmt_923: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_926_wire & type_cast_929_wire_constant;
      req <= phi_stmt_923_req_0 & phi_stmt_923_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_923_ack_0,
          idata => idata,
          odata => i3x_x0x_xlcssa53_923,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_923
    addr_of_768_final_reg: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_767_root_address, dout => tmp12_769, req => addr_of_768_final_reg_req_0, ack => addr_of_768_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_804_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_803_root_address, dout => tmp17_805, req => addr_of_804_final_reg_req_0, ack => addr_of_804_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_934_final_reg: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_933_root_address, dout => tmp38_935, req => addr_of_934_final_reg_req_0, ack => addr_of_934_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_767_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => iNsTr_12_741, dout => simple_obj_ref_766_resized, req => array_obj_ref_767_index_0_resize_req_0, ack => array_obj_ref_767_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_767_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_766_scaled, dout => array_obj_ref_767_final_offset, req => array_obj_ref_767_offset_inst_req_0, ack => array_obj_ref_767_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_803_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp16_800, dout => simple_obj_ref_802_resized, req => array_obj_ref_803_index_0_resize_req_0, ack => array_obj_ref_803_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_803_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_802_scaled, dout => array_obj_ref_803_final_offset, req => array_obj_ref_803_offset_inst_req_0, ack => array_obj_ref_803_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_933_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => i3x_x0x_xlcssa53_923, dout => simple_obj_ref_932_resized, req => array_obj_ref_933_index_0_resize_req_0, ack => array_obj_ref_933_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_933_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_932_scaled, dout => array_obj_ref_933_final_offset, req => array_obj_ref_933_offset_inst_req_0, ack => array_obj_ref_933_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_772_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp12_769, dout => ptr_deref_772_resized_base_address, req => ptr_deref_772_base_resize_req_0, ack => ptr_deref_772_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_811_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp12_769, dout => ptr_deref_811_resized_base_address, req => ptr_deref_811_base_resize_req_0, ack => ptr_deref_811_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_937_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp38_935, dout => ptr_deref_937_resized_base_address, req => ptr_deref_937_base_resize_req_0, ack => ptr_deref_937_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_744_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp21_792, dout => type_cast_744_wire, req => type_cast_744_inst_req_0, ack => type_cast_744_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_752_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_12_741, dout => type_cast_752_wire, req => type_cast_752_inst_req_0, ack => type_cast_752_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_808_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_805, dout => tmp18_809, req => type_cast_808_inst_req_0, ack => type_cast_808_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_873_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_20_889, dout => type_cast_873_wire, req => type_cast_873_inst_req_0, ack => type_cast_873_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_910_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_20_889, dout => type_cast_910_wire, req => type_cast_910_inst_req_0, ack => type_cast_910_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_926_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_20_889, dout => type_cast_926_wire, req => type_cast_926_inst_req_0, ack => type_cast_926_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_767_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_767_index_0_rename_ack_0 <= array_obj_ref_767_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_766_resized;
      simple_obj_ref_766_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_767_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_767_root_address_inst_ack_0 <= array_obj_ref_767_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_767_final_offset;
      array_obj_ref_767_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_803_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_803_index_0_rename_ack_0 <= array_obj_ref_803_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_802_resized;
      simple_obj_ref_802_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_933_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_933_index_0_rename_ack_0 <= array_obj_ref_933_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_932_resized;
      simple_obj_ref_932_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_933_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_933_root_address_inst_ack_0 <= array_obj_ref_933_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_933_final_offset;
      array_obj_ref_933_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_682_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_682_gather_scatter_ack_0 <= ptr_deref_682_gather_scatter_req_0;
      aggregated_sig <= type_cast_684_wire_constant;
      ptr_deref_682_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_693_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_693_gather_scatter_ack_0 <= ptr_deref_693_gather_scatter_req_0;
      aggregated_sig <= type_cast_695_wire_constant;
      ptr_deref_693_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_704_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_704_gather_scatter_ack_0 <= ptr_deref_704_gather_scatter_req_0;
      aggregated_sig <= type_cast_706_wire_constant;
      ptr_deref_704_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_715_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_715_gather_scatter_ack_0 <= ptr_deref_715_gather_scatter_req_0;
      aggregated_sig <= type_cast_717_wire_constant;
      ptr_deref_715_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_772_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_772_addr_0_ack_0 <= ptr_deref_772_addr_0_req_0;
      aggregated_sig <= ptr_deref_772_root_address;
      ptr_deref_772_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_772_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_772_gather_scatter_ack_0 <= ptr_deref_772_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_772_data_0;
      tmp13_773 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_772_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_772_root_address_inst_ack_0 <= ptr_deref_772_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_772_resized_base_address;
      ptr_deref_772_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_811_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_811_addr_0_ack_0 <= ptr_deref_811_addr_0_req_0;
      aggregated_sig <= ptr_deref_811_root_address;
      ptr_deref_811_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_811_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_811_gather_scatter_ack_0 <= ptr_deref_811_gather_scatter_req_0;
      aggregated_sig <= type_cast_813_wire_constant;
      ptr_deref_811_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_811_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_811_root_address_inst_ack_0 <= ptr_deref_811_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_811_resized_base_address;
      ptr_deref_811_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_937_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_937_addr_0_ack_0 <= ptr_deref_937_addr_0_req_0;
      aggregated_sig <= ptr_deref_937_root_address;
      ptr_deref_937_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_937_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_937_gather_scatter_ack_0 <= ptr_deref_937_gather_scatter_req_0;
      aggregated_sig <= type_cast_939_wire_constant;
      ptr_deref_937_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_937_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_937_root_address_inst_ack_0 <= ptr_deref_937_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_937_resized_base_address;
      ptr_deref_937_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    if_stmt_758_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp10_757;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_758_branch_req_0,
          ack0 => if_stmt_758_branch_ack_0,
          ack1 => if_stmt_758_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_780_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp14_779;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_780_branch_req_0,
          ack0 => if_stmt_780_branch_ack_0,
          ack1 => if_stmt_780_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_863_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp3243_862;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_863_branch_req_0,
          ack0 => if_stmt_863_branch_ack_0,
          ack1 => if_stmt_863_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_901_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp32_900;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_901_branch_req_0,
          ack0 => if_stmt_901_branch_ack_0,
          ack1 => if_stmt_901_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_916_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp36_915;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_916_branch_req_0,
          ack0 => if_stmt_916_branch_ack_0,
          ack1 => if_stmt_916_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_730_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_732_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_730_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_730_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_730_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_735_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_730_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_730_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_730_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_732_wire_constant_cmp & expr_735_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_730_branch_default_req_0,
          ack0 => switch_stmt_730_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_803_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_803_final_offset;
      array_obj_ref_803_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_803_root_address_inst_req_0,
          ackL => array_obj_ref_803_root_address_inst_ack_0,
          reqR => array_obj_ref_803_root_address_inst_req_1,
          ackR => array_obj_ref_803_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_756_inst binary_914_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_752_wire & type_cast_910_wire;
      tmp10_757 <= data_out(1 downto 1);
      tmp36_915 <= data_out(0 downto 0);
      reqL(1) <= binary_756_inst_req_0;
      reqL(0) <= binary_914_inst_req_0;
      binary_756_inst_ack_0 <= ackL(1);
      binary_914_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_756_inst_req_1;
      reqR(0) <= binary_914_inst_req_1;
      binary_756_inst_ack_1 <= ackR(1);
      binary_914_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : switch_stmt_730_select_expr_1 binary_778_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_729 & tmp13_773;
      expr_735_wire_constant_cmp <= data_out(1 downto 1);
      tmp14_779 <= data_out(0 downto 0);
      reqL(1) <= switch_stmt_730_select_expr_1_req_0;
      reqL(0) <= binary_778_inst_req_0;
      switch_stmt_730_select_expr_1_ack_0 <= ackL(1);
      binary_778_inst_ack_0 <= ackL(0);
      reqR(1) <= switch_stmt_730_select_expr_1_req_1;
      reqR(0) <= binary_778_inst_req_1;
      switch_stmt_730_select_expr_1_ack_1 <= ackR(1);
      binary_778_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_888_inst binary_791_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= i3x_x044_870 & iNsTr_12_741;
      iNsTr_20_889 <= data_out(63 downto 32);
      tmp21_792 <= data_out(31 downto 0);
      reqL(1) <= binary_888_inst_req_0;
      reqL(0) <= binary_791_inst_req_0;
      binary_888_inst_ack_0 <= ackL(1);
      binary_791_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_888_inst_req_1;
      reqR(0) <= binary_791_inst_req_1;
      binary_888_inst_ack_1 <= ackR(1);
      binary_791_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_799_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_741;
      tmp16_800 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_799_inst_req_0,
          ackL => binary_799_inst_ack_0,
          reqR => binary_799_inst_req_1,
          ackR => binary_799_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_861_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp28_856;
      tmp3243_862 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000100000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_861_inst_req_0,
          ackL => binary_861_inst_ack_0,
          reqR => binary_861_inst_req_1,
          ackR => binary_861_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_882_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= i3x_x044_870;
      tmp50_883 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_882_inst_req_0,
          ackL => binary_882_inst_ack_0,
          reqR => binary_882_inst_req_1,
          ackR => binary_882_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_894_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp50_883;
      tmp31_895 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000001000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_894_inst_req_0,
          ackL => binary_894_inst_ack_0,
          reqR => binary_894_inst_req_1,
          ackR => binary_894_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_899_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp28_856 & tmp31_895;
      tmp32_900 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_899_inst_req_0,
          ackL => binary_899_inst_ack_0,
          reqR => binary_899_inst_req_1,
          ackR => binary_899_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : switch_stmt_730_select_expr_0 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_729;
      expr_732_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000010",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_730_select_expr_0_req_0,
          ackL => switch_stmt_730_select_expr_0_ack_0,
          reqR => switch_stmt_730_select_expr_0_req_1,
          ackR => switch_stmt_730_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared load operator group (0) : ptr_deref_772_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_772_load_0_req_0;
      ptr_deref_772_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_772_load_0_req_1;
      ptr_deref_772_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_772_word_address_0;
      ptr_deref_772_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 3,  num_reqs => 1,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(2 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_682_store_0 ptr_deref_811_store_0 ptr_deref_937_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(8 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_682_store_0_req_0;
      reqL(1) <= ptr_deref_811_store_0_req_0;
      reqL(0) <= ptr_deref_937_store_0_req_0;
      ptr_deref_682_store_0_ack_0 <= ackL(2);
      ptr_deref_811_store_0_ack_0 <= ackL(1);
      ptr_deref_937_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_682_store_0_req_1;
      reqR(1) <= ptr_deref_811_store_0_req_1;
      reqR(0) <= ptr_deref_937_store_0_req_1;
      ptr_deref_682_store_0_ack_1 <= ackR(2);
      ptr_deref_811_store_0_ack_1 <= ackR(1);
      ptr_deref_937_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_682_word_address_0 & ptr_deref_811_word_address_0 & ptr_deref_937_word_address_0;
      data_in <= ptr_deref_682_data_0 & ptr_deref_811_data_0 & ptr_deref_937_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(3),
          mack => memory_space_2_sr_ack(3),
          maddr => memory_space_2_sr_addr(11 downto 9),
          mdata => memory_space_2_sr_data(31 downto 24),
          mtag => memory_space_2_sr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(3),
          mack => memory_space_2_sc_ack(3),
          mtag => memory_space_2_sc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_693_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_693_store_0_req_0;
      ptr_deref_693_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_693_store_0_req_1;
      ptr_deref_693_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_693_word_address_0;
      data_in <= ptr_deref_693_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(2),
          mack => memory_space_2_sr_ack(2),
          maddr => memory_space_2_sr_addr(8 downto 6),
          mdata => memory_space_2_sr_data(23 downto 16),
          mtag => memory_space_2_sr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(2),
          mack => memory_space_2_sc_ack(2),
          mtag => memory_space_2_sc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_704_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_704_store_0_req_0;
      ptr_deref_704_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_704_store_0_req_1;
      ptr_deref_704_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_704_word_address_0;
      data_in <= ptr_deref_704_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(1),
          mack => memory_space_2_sr_ack(1),
          maddr => memory_space_2_sr_addr(5 downto 3),
          mdata => memory_space_2_sr_data(15 downto 8),
          mtag => memory_space_2_sr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(1),
          mack => memory_space_2_sc_ack(1),
          mtag => memory_space_2_sc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_715_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_715_store_0_req_0;
      ptr_deref_715_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_715_store_0_req_1;
      ptr_deref_715_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_715_word_address_0;
      data_in <= ptr_deref_715_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(2 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : simple_obj_ref_728_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_728_inst_req_0;
      simple_obj_ref_728_inst_ack_0 <= ack(0);
      tmp6_729 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_request_pipe_read_req(0),
          oack => free_queue_request_pipe_read_ack(0),
          odata => free_queue_request_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_855_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_855_inst_req_0;
      simple_obj_ref_855_inst_ack_0 <= ack(0);
      tmp28_856 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_put_pipe_read_req(0),
          oack => free_queue_put_pipe_read_ack(0),
          odata => free_queue_put_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_821_inst simple_obj_ref_842_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_821_inst_req_0;
      req(0) <= simple_obj_ref_842_inst_req_0;
      simple_obj_ref_821_inst_ack_0 <= ack(1);
      simple_obj_ref_842_inst_ack_0 <= ack(0);
      data_in <= type_cast_823_wire_constant & type_cast_844_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 2,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_ack_pipe_write_req(0),
          oack => free_queue_ack_pipe_write_ack(0),
          odata => free_queue_ack_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_831_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_831_inst_req_0;
      simple_obj_ref_831_inst_ack_0 <= ack(0);
      data_in <= tmp18_809;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_get_pipe_write_req(0),
          oack => free_queue_get_pipe_write_ack(0),
          odata => free_queue_get_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_674_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_674_call_req_0;
      call_stmt_674_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_674_call_req_1;
      call_stmt_674_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => global_storage_initializer_x_call_reqs(0),
          ackR => global_storage_initializer_x_call_acks(0),
          tagR => global_storage_initializer_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => global_storage_initializer_x_return_acks(0), -- cross-over
          ackL => global_storage_initializer_x_return_reqs(0), -- cross-over
          tagL => global_storage_initializer_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity global_storage_initializer_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    default_initializer_xx_xstr2_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr2_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr4_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_foo_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_foo_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_foo_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_foo_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_foo_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_foo_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_free_queue_ram_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr5_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr8_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr7_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr1_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr3_return_tag :  in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_call_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_call_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_call_tag  :  out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_return_reqs : out  std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_return_acks : in   std_logic_vector(0 downto 0);
    default_initializer_xx_xstr6_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity global_storage_initializer_x;
architecture Default of global_storage_initializer_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal global_storage_initializer_x_xCP_2874_start: Boolean;
  -- links between control-path and data-path
  signal call_stmt_946_call_req_0 : boolean;
  signal call_stmt_946_call_ack_0 : boolean;
  signal call_stmt_946_call_req_1 : boolean;
  signal call_stmt_946_call_ack_1 : boolean;
  signal call_stmt_947_call_req_0 : boolean;
  signal call_stmt_947_call_ack_0 : boolean;
  signal call_stmt_947_call_req_1 : boolean;
  signal call_stmt_947_call_ack_1 : boolean;
  signal call_stmt_948_call_req_0 : boolean;
  signal call_stmt_948_call_ack_0 : boolean;
  signal call_stmt_948_call_req_1 : boolean;
  signal call_stmt_948_call_ack_1 : boolean;
  signal call_stmt_949_call_req_0 : boolean;
  signal call_stmt_949_call_ack_0 : boolean;
  signal call_stmt_949_call_req_1 : boolean;
  signal call_stmt_949_call_ack_1 : boolean;
  signal call_stmt_950_call_req_0 : boolean;
  signal call_stmt_950_call_ack_0 : boolean;
  signal call_stmt_950_call_req_1 : boolean;
  signal call_stmt_950_call_ack_1 : boolean;
  signal call_stmt_951_call_req_0 : boolean;
  signal call_stmt_951_call_ack_0 : boolean;
  signal call_stmt_951_call_req_1 : boolean;
  signal call_stmt_951_call_ack_1 : boolean;
  signal call_stmt_952_call_req_0 : boolean;
  signal call_stmt_952_call_ack_0 : boolean;
  signal call_stmt_952_call_req_1 : boolean;
  signal call_stmt_952_call_ack_1 : boolean;
  signal call_stmt_953_call_req_0 : boolean;
  signal call_stmt_953_call_ack_0 : boolean;
  signal call_stmt_953_call_req_1 : boolean;
  signal call_stmt_953_call_ack_1 : boolean;
  signal call_stmt_954_call_req_0 : boolean;
  signal call_stmt_954_call_ack_0 : boolean;
  signal call_stmt_954_call_req_1 : boolean;
  signal call_stmt_954_call_ack_1 : boolean;
  signal call_stmt_955_call_req_0 : boolean;
  signal call_stmt_955_call_ack_0 : boolean;
  signal call_stmt_955_call_req_1 : boolean;
  signal call_stmt_955_call_ack_1 : boolean;
  signal call_stmt_956_call_req_0 : boolean;
  signal call_stmt_956_call_ack_0 : boolean;
  signal call_stmt_956_call_req_1 : boolean;
  signal call_stmt_956_call_ack_1 : boolean;
  signal call_stmt_957_call_req_0 : boolean;
  signal call_stmt_957_call_ack_0 : boolean;
  signal call_stmt_957_call_req_1 : boolean;
  signal call_stmt_957_call_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  global_storage_initializer_x_xCP_2874: Block -- control-path 
    signal cp_elements: BooleanArray(37 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(37);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(37), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    call_stmt_946_call_req_0 <= cp_elements(1);
    cp_elements(2) <= call_stmt_946_call_ack_0;
    call_stmt_946_call_req_1 <= cp_elements(2);
    cp_elements(3) <= call_stmt_946_call_ack_1;
    cp_elements(4) <= cp_elements(0);
    call_stmt_947_call_req_0 <= cp_elements(4);
    cp_elements(5) <= call_stmt_947_call_ack_0;
    call_stmt_947_call_req_1 <= cp_elements(5);
    cp_elements(6) <= call_stmt_947_call_ack_1;
    cp_elements(7) <= cp_elements(0);
    call_stmt_948_call_req_0 <= cp_elements(7);
    cp_elements(8) <= call_stmt_948_call_ack_0;
    call_stmt_948_call_req_1 <= cp_elements(8);
    cp_elements(9) <= call_stmt_948_call_ack_1;
    cp_elements(10) <= cp_elements(0);
    call_stmt_949_call_req_0 <= cp_elements(10);
    cp_elements(11) <= call_stmt_949_call_ack_0;
    call_stmt_949_call_req_1 <= cp_elements(11);
    cp_elements(12) <= call_stmt_949_call_ack_1;
    cp_elements(13) <= cp_elements(0);
    call_stmt_950_call_req_0 <= cp_elements(13);
    cp_elements(14) <= call_stmt_950_call_ack_0;
    call_stmt_950_call_req_1 <= cp_elements(14);
    cp_elements(15) <= call_stmt_950_call_ack_1;
    cp_elements(16) <= cp_elements(0);
    call_stmt_951_call_req_0 <= cp_elements(16);
    cp_elements(17) <= call_stmt_951_call_ack_0;
    call_stmt_951_call_req_1 <= cp_elements(17);
    cp_elements(18) <= call_stmt_951_call_ack_1;
    cp_elements(19) <= cp_elements(0);
    call_stmt_952_call_req_0 <= cp_elements(19);
    cp_elements(20) <= call_stmt_952_call_ack_0;
    call_stmt_952_call_req_1 <= cp_elements(20);
    cp_elements(21) <= call_stmt_952_call_ack_1;
    cp_elements(22) <= cp_elements(0);
    call_stmt_953_call_req_0 <= cp_elements(22);
    cp_elements(23) <= call_stmt_953_call_ack_0;
    call_stmt_953_call_req_1 <= cp_elements(23);
    cp_elements(24) <= call_stmt_953_call_ack_1;
    cp_elements(25) <= cp_elements(0);
    call_stmt_954_call_req_0 <= cp_elements(25);
    cp_elements(26) <= call_stmt_954_call_ack_0;
    call_stmt_954_call_req_1 <= cp_elements(26);
    cp_elements(27) <= call_stmt_954_call_ack_1;
    cp_elements(28) <= cp_elements(0);
    call_stmt_955_call_req_0 <= cp_elements(28);
    cp_elements(29) <= call_stmt_955_call_ack_0;
    call_stmt_955_call_req_1 <= cp_elements(29);
    cp_elements(30) <= call_stmt_955_call_ack_1;
    cp_elements(31) <= cp_elements(0);
    call_stmt_956_call_req_0 <= cp_elements(31);
    cp_elements(32) <= call_stmt_956_call_ack_0;
    call_stmt_956_call_req_1 <= cp_elements(32);
    cp_elements(33) <= call_stmt_956_call_ack_1;
    cp_elements(34) <= cp_elements(0);
    call_stmt_957_call_req_0 <= cp_elements(34);
    cp_elements(35) <= call_stmt_957_call_ack_0;
    call_stmt_957_call_req_1 <= cp_elements(35);
    cp_elements(36) <= call_stmt_957_call_ack_1;
    cpelement_group_37 : Block -- 
      signal predecessors: BooleanArray(11 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(6) & cp_elements(9) & cp_elements(12) & cp_elements(15) & cp_elements(18) & cp_elements(21) & cp_elements(24) & cp_elements(27) & cp_elements(30) & cp_elements(33) & cp_elements(36));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(37),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared call operator group (0) : call_stmt_946_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_946_call_req_0;
      call_stmt_946_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_946_call_req_1;
      call_stmt_946_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr_call_reqs(0),
          ackR => default_initializer_xx_xstr_call_acks(0),
          tagR => default_initializer_xx_xstr_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_947_call 
    CallGroup1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_947_call_req_0;
      call_stmt_947_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_947_call_req_1;
      call_stmt_947_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr1_call_reqs(0),
          ackR => default_initializer_xx_xstr1_call_acks(0),
          tagR => default_initializer_xx_xstr1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr1_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr1_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_948_call 
    CallGroup2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_948_call_req_0;
      call_stmt_948_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_948_call_req_1;
      call_stmt_948_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr2_call_reqs(0),
          ackR => default_initializer_xx_xstr2_call_acks(0),
          tagR => default_initializer_xx_xstr2_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr2_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr2_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr2_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_949_call 
    CallGroup3: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_949_call_req_0;
      call_stmt_949_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_949_call_req_1;
      call_stmt_949_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr3_call_reqs(0),
          ackR => default_initializer_xx_xstr3_call_acks(0),
          tagR => default_initializer_xx_xstr3_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr3_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr3_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr3_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_950_call 
    CallGroup4: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_950_call_req_0;
      call_stmt_950_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_950_call_req_1;
      call_stmt_950_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_free_queue_call_reqs(0),
          ackR => default_initializer_free_queue_call_acks(0),
          tagR => default_initializer_free_queue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_free_queue_return_acks(0), -- cross-over
          ackL => default_initializer_free_queue_return_reqs(0), -- cross-over
          tagL => default_initializer_free_queue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_951_call 
    CallGroup5: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_951_call_req_0;
      call_stmt_951_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_951_call_req_1;
      call_stmt_951_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_free_queue_ram_call_reqs(0),
          ackR => default_initializer_free_queue_ram_call_acks(0),
          tagR => default_initializer_free_queue_ram_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_free_queue_ram_return_acks(0), -- cross-over
          ackL => default_initializer_free_queue_ram_return_reqs(0), -- cross-over
          tagL => default_initializer_free_queue_ram_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_952_call 
    CallGroup6: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_952_call_req_0;
      call_stmt_952_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_952_call_req_1;
      call_stmt_952_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_foo_call_reqs(0),
          ackR => default_initializer_foo_call_acks(0),
          tagR => default_initializer_foo_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_foo_return_acks(0), -- cross-over
          ackL => default_initializer_foo_return_reqs(0), -- cross-over
          tagL => default_initializer_foo_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_953_call 
    CallGroup7: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_953_call_req_0;
      call_stmt_953_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_953_call_req_1;
      call_stmt_953_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr4_call_reqs(0),
          ackR => default_initializer_xx_xstr4_call_acks(0),
          tagR => default_initializer_xx_xstr4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr4_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr4_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_954_call 
    CallGroup8: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_954_call_req_0;
      call_stmt_954_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_954_call_req_1;
      call_stmt_954_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr5_call_reqs(0),
          ackR => default_initializer_xx_xstr5_call_acks(0),
          tagR => default_initializer_xx_xstr5_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr5_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr5_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr5_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- shared call operator group (9) : call_stmt_955_call 
    CallGroup9: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_955_call_req_0;
      call_stmt_955_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_955_call_req_1;
      call_stmt_955_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr6_call_reqs(0),
          ackR => default_initializer_xx_xstr6_call_acks(0),
          tagR => default_initializer_xx_xstr6_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr6_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr6_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr6_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 9
    -- shared call operator group (10) : call_stmt_956_call 
    CallGroup10: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_956_call_req_0;
      call_stmt_956_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_956_call_req_1;
      call_stmt_956_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr7_call_reqs(0),
          ackR => default_initializer_xx_xstr7_call_acks(0),
          tagR => default_initializer_xx_xstr7_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr7_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr7_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr7_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 10
    -- shared call operator group (11) : call_stmt_957_call 
    CallGroup11: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_957_call_req_0;
      call_stmt_957_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_957_call_req_1;
      call_stmt_957_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => default_initializer_xx_xstr8_call_reqs(0),
          ackR => default_initializer_xx_xstr8_call_acks(0),
          tagR => default_initializer_xx_xstr8_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => default_initializer_xx_xstr8_return_acks(0), -- cross-over
          ackL => default_initializer_xx_xstr8_return_reqs(0), -- cross-over
          tagL => default_initializer_xx_xstr8_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 11
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_input is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_0_sr_req : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(7 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(87 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(15 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(7 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(7 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(15 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
    in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    midpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    midpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    midpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_input;
architecture Default of wrapper_input is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_input_CP_4300_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_969_store_0_ack_0 : boolean;
  signal ptr_deref_1231_store_0_ack_0 : boolean;
  signal ptr_deref_1245_store_0_req_0 : boolean;
  signal ptr_deref_1281_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1014_inst_ack_0 : boolean;
  signal ptr_deref_969_store_0_req_0 : boolean;
  signal binary_1266_inst_ack_0 : boolean;
  signal ptr_deref_1245_store_0_ack_0 : boolean;
  signal ptr_deref_1245_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1259_store_0_ack_1 : boolean;
  signal type_cast_1023_inst_ack_0 : boolean;
  signal type_cast_1256_inst_req_0 : boolean;
  signal type_cast_1256_inst_ack_0 : boolean;
  signal simple_obj_ref_1014_inst_req_0 : boolean;
  signal ptr_deref_1217_base_resize_ack_0 : boolean;
  signal simple_obj_ref_981_inst_ack_0 : boolean;
  signal binary_998_inst_req_1 : boolean;
  signal ptr_deref_1217_base_resize_req_0 : boolean;
  signal binary_1266_inst_req_1 : boolean;
  signal array_obj_ref_1043_base_resize_req_0 : boolean;
  signal array_obj_ref_1048_base_resize_ack_0 : boolean;
  signal ptr_deref_1281_addr_0_ack_0 : boolean;
  signal ptr_deref_1245_addr_0_ack_0 : boolean;
  signal ptr_deref_1259_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_992_inst_ack_0 : boolean;
  signal ptr_deref_1259_addr_0_ack_0 : boolean;
  signal array_obj_ref_1033_root_address_inst_ack_1 : boolean;
  signal binary_1418_inst_req_0 : boolean;
  signal array_obj_ref_1028_final_reg_ack_0 : boolean;
  signal binary_998_inst_req_0 : boolean;
  signal array_obj_ref_1038_base_resize_ack_0 : boolean;
  signal ptr_deref_1231_addr_0_req_0 : boolean;
  signal simple_obj_ref_981_inst_req_0 : boolean;
  signal array_obj_ref_1033_base_resize_ack_0 : boolean;
  signal ptr_deref_1259_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1028_base_resize_req_0 : boolean;
  signal type_cast_1228_inst_ack_0 : boolean;
  signal if_stmt_1000_branch_req_0 : boolean;
  signal array_obj_ref_1048_final_reg_ack_0 : boolean;
  signal ptr_deref_1281_root_address_inst_ack_0 : boolean;
  signal type_cast_1278_inst_ack_0 : boolean;
  signal type_cast_1023_inst_req_0 : boolean;
  signal ptr_deref_1217_addr_0_req_0 : boolean;
  signal ptr_deref_1245_addr_0_req_0 : boolean;
  signal array_obj_ref_1446_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1245_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1245_store_0_ack_1 : boolean;
  signal ptr_deref_1231_store_0_req_0 : boolean;
  signal binary_1266_inst_req_0 : boolean;
  signal array_obj_ref_1033_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1048_final_reg_req_0 : boolean;
  signal binary_1224_inst_req_1 : boolean;
  signal binary_1224_inst_ack_0 : boolean;
  signal array_obj_ref_1028_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1217_addr_0_ack_0 : boolean;
  signal ptr_deref_1259_base_resize_ack_0 : boolean;
  signal ptr_deref_1259_addr_0_req_0 : boolean;
  signal ptr_deref_1425_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1273_store_0_ack_0 : boolean;
  signal ptr_deref_1231_addr_0_ack_0 : boolean;
  signal binary_998_inst_ack_0 : boolean;
  signal array_obj_ref_1043_final_reg_ack_0 : boolean;
  signal ptr_deref_1231_base_resize_req_0 : boolean;
  signal ptr_deref_969_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1281_base_resize_ack_0 : boolean;
  signal ptr_deref_1259_store_0_ack_0 : boolean;
  signal array_obj_ref_1038_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1449_gather_scatter_ack_0 : boolean;
  signal type_cast_1270_inst_req_0 : boolean;
  signal array_obj_ref_1033_base_resize_req_0 : boolean;
  signal binary_1266_inst_ack_1 : boolean;
  signal ptr_deref_969_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1028_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1033_root_address_inst_req_1 : boolean;
  signal binary_998_inst_ack_1 : boolean;
  signal ptr_deref_1231_base_resize_ack_0 : boolean;
  signal type_cast_1242_inst_ack_0 : boolean;
  signal ptr_deref_1273_store_0_req_0 : boolean;
  signal ptr_deref_1281_store_0_ack_0 : boolean;
  signal ptr_deref_1245_base_resize_ack_0 : boolean;
  signal binary_1290_inst_req_0 : boolean;
  signal ptr_deref_1281_base_resize_req_0 : boolean;
  signal type_cast_1018_inst_req_0 : boolean;
  signal ptr_deref_1259_base_resize_req_0 : boolean;
  signal ptr_deref_1259_store_0_req_1 : boolean;
  signal type_cast_1052_inst_req_0 : boolean;
  signal type_cast_1242_inst_req_0 : boolean;
  signal type_cast_1270_inst_ack_0 : boolean;
  signal array_obj_ref_1048_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1245_store_0_req_1 : boolean;
  signal binary_1224_inst_ack_1 : boolean;
  signal array_obj_ref_1048_root_address_inst_req_1 : boolean;
  signal ptr_deref_1217_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1043_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1057_base_resize_ack_0 : boolean;
  signal ptr_deref_1281_store_0_req_1 : boolean;
  signal binary_1418_inst_req_1 : boolean;
  signal type_cast_1018_inst_ack_0 : boolean;
  signal array_obj_ref_1048_root_address_inst_ack_1 : boolean;
  signal type_cast_1228_inst_req_0 : boolean;
  signal ptr_deref_1425_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1043_root_address_inst_ack_0 : boolean;
  signal binary_1466_inst_ack_1 : boolean;
  signal ptr_deref_1273_store_0_ack_1 : boolean;
  signal array_obj_ref_1043_final_reg_req_0 : boolean;
  signal array_obj_ref_1038_root_address_inst_req_1 : boolean;
  signal ptr_deref_969_store_0_req_1 : boolean;
  signal ptr_deref_1381_root_address_inst_req_0 : boolean;
  signal ptr_deref_1425_addr_0_req_0 : boolean;
  signal type_cast_1278_inst_req_0 : boolean;
  signal ptr_deref_969_store_0_ack_1 : boolean;
  signal if_stmt_1000_branch_ack_1 : boolean;
  signal array_obj_ref_1028_root_address_inst_req_0 : boolean;
  signal binary_1418_inst_ack_1 : boolean;
  signal array_obj_ref_1038_final_reg_req_0 : boolean;
  signal array_obj_ref_1048_base_resize_req_0 : boolean;
  signal ptr_deref_1273_store_0_req_1 : boolean;
  signal ptr_deref_1259_root_address_inst_ack_0 : boolean;
  signal if_stmt_1000_branch_ack_0 : boolean;
  signal array_obj_ref_1043_base_resize_ack_0 : boolean;
  signal ptr_deref_1389_store_0_ack_1 : boolean;
  signal ptr_deref_1281_store_0_req_0 : boolean;
  signal array_obj_ref_1028_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1033_final_reg_req_0 : boolean;
  signal ptr_deref_1231_root_address_inst_req_0 : boolean;
  signal binary_1252_inst_ack_1 : boolean;
  signal array_obj_ref_1038_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1259_store_0_req_0 : boolean;
  signal ptr_deref_1245_root_address_inst_req_0 : boolean;
  signal binary_1252_inst_req_1 : boolean;
  signal ptr_deref_1245_gather_scatter_req_0 : boolean;
  signal ptr_deref_1245_base_resize_req_0 : boolean;
  signal ptr_deref_1217_store_0_ack_0 : boolean;
  signal binary_1252_inst_ack_0 : boolean;
  signal ptr_deref_1259_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1038_base_resize_req_0 : boolean;
  signal array_obj_ref_1028_base_resize_ack_0 : boolean;
  signal array_obj_ref_1033_final_reg_ack_0 : boolean;
  signal ptr_deref_1449_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1038_final_reg_ack_0 : boolean;
  signal ptr_deref_1231_gather_scatter_ack_0 : boolean;
  signal binary_1252_inst_req_0 : boolean;
  signal ptr_deref_1231_gather_scatter_req_0 : boolean;
  signal ptr_deref_1381_base_resize_ack_0 : boolean;
  signal type_cast_1052_inst_ack_0 : boolean;
  signal array_obj_ref_1033_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1470_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1217_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1281_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_992_inst_req_0 : boolean;
  signal array_obj_ref_1048_root_address_inst_req_0 : boolean;
  signal ptr_deref_1273_gather_scatter_ack_0 : boolean;
  signal binary_1238_inst_ack_0 : boolean;
  signal ptr_deref_1273_gather_scatter_req_0 : boolean;
  signal binary_1238_inst_req_0 : boolean;
  signal binary_1238_inst_ack_1 : boolean;
  signal binary_1238_inst_req_1 : boolean;
  signal ptr_deref_1389_store_0_req_1 : boolean;
  signal array_obj_ref_1470_base_resize_req_0 : boolean;
  signal ptr_deref_1425_addr_0_ack_0 : boolean;
  signal array_obj_ref_1062_final_reg_req_0 : boolean;
  signal ptr_deref_1273_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1062_final_reg_ack_0 : boolean;
  signal binary_1290_inst_ack_1 : boolean;
  signal array_obj_ref_1067_final_reg_req_0 : boolean;
  signal array_obj_ref_1067_final_reg_ack_0 : boolean;
  signal array_obj_ref_1067_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1067_root_address_inst_ack_1 : boolean;
  signal type_cast_1294_inst_req_0 : boolean;
  signal array_obj_ref_1057_base_resize_req_0 : boolean;
  signal ptr_deref_1231_store_0_ack_1 : boolean;
  signal array_obj_ref_1446_base_resize_req_0 : boolean;
  signal array_obj_ref_1067_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1067_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1231_store_0_req_1 : boolean;
  signal binary_1466_inst_ack_0 : boolean;
  signal array_obj_ref_1057_root_address_inst_req_1 : boolean;
  signal type_cast_1214_inst_req_0 : boolean;
  signal array_obj_ref_1057_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1470_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1281_root_address_inst_req_0 : boolean;
  signal ptr_deref_1273_base_resize_ack_0 : boolean;
  signal ptr_deref_1273_base_resize_req_0 : boolean;
  signal array_obj_ref_1057_final_reg_req_0 : boolean;
  signal ptr_deref_1389_base_resize_req_0 : boolean;
  signal ptr_deref_1381_addr_0_ack_0 : boolean;
  signal ptr_deref_1273_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1470_final_reg_ack_0 : boolean;
  signal ptr_deref_1217_store_0_req_1 : boolean;
  signal ptr_deref_1273_addr_0_ack_0 : boolean;
  signal array_obj_ref_1062_root_address_inst_req_0 : boolean;
  signal ptr_deref_1273_addr_0_req_0 : boolean;
  signal array_obj_ref_1062_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1062_root_address_inst_req_1 : boolean;
  signal ptr_deref_1217_store_0_ack_1 : boolean;
  signal array_obj_ref_1062_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1470_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1062_base_resize_req_0 : boolean;
  signal array_obj_ref_1062_base_resize_ack_0 : boolean;
  signal ptr_deref_1425_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1057_final_reg_ack_0 : boolean;
  signal ptr_deref_1381_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1043_root_address_inst_ack_1 : boolean;
  signal type_cast_1214_inst_ack_0 : boolean;
  signal array_obj_ref_1043_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1446_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1057_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1057_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1067_base_resize_req_0 : boolean;
  signal array_obj_ref_1067_base_resize_ack_0 : boolean;
  signal ptr_deref_1381_base_resize_req_0 : boolean;
  signal binary_1224_inst_req_0 : boolean;
  signal array_obj_ref_1038_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1028_final_reg_req_0 : boolean;
  signal ptr_deref_1231_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1217_gather_scatter_req_0 : boolean;
  signal binary_1290_inst_req_1 : boolean;
  signal ptr_deref_1217_gather_scatter_ack_0 : boolean;
  signal binary_1290_inst_ack_0 : boolean;
  signal ptr_deref_1425_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1281_store_0_ack_1 : boolean;
  signal ptr_deref_1281_addr_0_req_0 : boolean;
  signal ptr_deref_1217_store_0_req_0 : boolean;
  signal type_cast_1460_inst_ack_0 : boolean;
  signal binary_1466_inst_req_0 : boolean;
  signal ptr_deref_1389_base_resize_ack_0 : boolean;
  signal binary_1083_inst_req_0 : boolean;
  signal binary_1083_inst_ack_0 : boolean;
  signal binary_1083_inst_req_1 : boolean;
  signal binary_1083_inst_ack_1 : boolean;
  signal binary_1089_inst_req_0 : boolean;
  signal binary_1089_inst_ack_0 : boolean;
  signal binary_1089_inst_req_1 : boolean;
  signal binary_1089_inst_ack_1 : boolean;
  signal ptr_deref_1381_addr_0_req_0 : boolean;
  signal ptr_deref_1425_store_0_req_0 : boolean;
  signal ptr_deref_1425_store_0_ack_0 : boolean;
  signal array_obj_ref_1446_base_resize_ack_0 : boolean;
  signal binary_1396_inst_req_0 : boolean;
  signal array_obj_ref_1093_index_0_resize_req_0 : boolean;
  signal ptr_deref_1449_store_0_req_0 : boolean;
  signal array_obj_ref_1093_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1093_index_0_scale_req_0 : boolean;
  signal binary_1396_inst_ack_0 : boolean;
  signal array_obj_ref_1093_index_0_scale_ack_0 : boolean;
  signal ptr_deref_1425_store_0_req_1 : boolean;
  signal array_obj_ref_1093_index_0_scale_req_1 : boolean;
  signal ptr_deref_1381_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1093_index_0_scale_ack_1 : boolean;
  signal binary_1396_inst_req_1 : boolean;
  signal array_obj_ref_1093_offset_inst_req_0 : boolean;
  signal array_obj_ref_1093_offset_inst_ack_0 : boolean;
  signal ptr_deref_1425_store_0_ack_1 : boolean;
  signal array_obj_ref_1093_base_resize_req_0 : boolean;
  signal array_obj_ref_1093_base_resize_ack_0 : boolean;
  signal ptr_deref_1381_gather_scatter_ack_0 : boolean;
  signal binary_1396_inst_ack_1 : boolean;
  signal ptr_deref_1449_store_0_ack_0 : boolean;
  signal array_obj_ref_1093_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1093_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1093_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1093_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1473_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1093_final_reg_req_0 : boolean;
  signal array_obj_ref_1093_final_reg_ack_0 : boolean;
  signal type_cast_1097_inst_req_0 : boolean;
  signal type_cast_1097_inst_ack_0 : boolean;
  signal array_obj_ref_1102_base_resize_req_0 : boolean;
  signal binary_1432_inst_req_0 : boolean;
  signal array_obj_ref_1102_base_resize_ack_0 : boolean;
  signal binary_1432_inst_ack_0 : boolean;
  signal binary_1432_inst_req_1 : boolean;
  signal binary_1432_inst_ack_1 : boolean;
  signal array_obj_ref_1102_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1102_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1102_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1102_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1102_final_reg_req_0 : boolean;
  signal array_obj_ref_1102_final_reg_ack_0 : boolean;
  signal type_cast_1402_inst_req_0 : boolean;
  signal type_cast_1402_inst_ack_0 : boolean;
  signal array_obj_ref_1107_base_resize_req_0 : boolean;
  signal array_obj_ref_1107_base_resize_ack_0 : boolean;
  signal array_obj_ref_1107_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1107_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1107_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1107_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1107_final_reg_req_0 : boolean;
  signal type_cast_1436_inst_req_0 : boolean;
  signal array_obj_ref_1107_final_reg_ack_0 : boolean;
  signal ptr_deref_1381_store_0_req_0 : boolean;
  signal type_cast_1436_inst_ack_0 : boolean;
  signal ptr_deref_1381_store_0_ack_0 : boolean;
  signal binary_1418_inst_ack_0 : boolean;
  signal array_obj_ref_1112_base_resize_req_0 : boolean;
  signal array_obj_ref_1112_base_resize_ack_0 : boolean;
  signal array_obj_ref_1112_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1112_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1449_store_0_req_1 : boolean;
  signal array_obj_ref_1112_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1112_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1473_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1112_final_reg_req_0 : boolean;
  signal array_obj_ref_1112_final_reg_ack_0 : boolean;
  signal array_obj_ref_1470_base_resize_ack_0 : boolean;
  signal binary_1408_inst_req_0 : boolean;
  signal ptr_deref_1449_store_0_ack_1 : boolean;
  signal binary_1408_inst_ack_0 : boolean;
  signal binary_1118_inst_req_0 : boolean;
  signal binary_1118_inst_ack_0 : boolean;
  signal binary_1118_inst_req_1 : boolean;
  signal binary_1118_inst_ack_1 : boolean;
  signal binary_1442_inst_req_0 : boolean;
  signal binary_1442_inst_ack_0 : boolean;
  signal binary_1442_inst_req_1 : boolean;
  signal binary_1442_inst_ack_1 : boolean;
  signal array_obj_ref_1122_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1122_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1122_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1122_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1122_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1122_index_0_scale_ack_1 : boolean;
  signal binary_1408_inst_req_1 : boolean;
  signal array_obj_ref_1470_final_reg_req_0 : boolean;
  signal array_obj_ref_1122_offset_inst_req_0 : boolean;
  signal array_obj_ref_1122_offset_inst_ack_0 : boolean;
  signal binary_1408_inst_ack_1 : boolean;
  signal array_obj_ref_1122_base_resize_req_0 : boolean;
  signal array_obj_ref_1122_base_resize_ack_0 : boolean;
  signal ptr_deref_1473_addr_0_req_0 : boolean;
  signal array_obj_ref_1122_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1122_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1122_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1122_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1381_store_0_req_1 : boolean;
  signal ptr_deref_1381_store_0_ack_1 : boolean;
  signal array_obj_ref_1122_final_reg_req_0 : boolean;
  signal array_obj_ref_1122_final_reg_ack_0 : boolean;
  signal type_cast_1126_inst_req_0 : boolean;
  signal type_cast_1126_inst_ack_0 : boolean;
  signal array_obj_ref_1131_base_resize_req_0 : boolean;
  signal array_obj_ref_1131_base_resize_ack_0 : boolean;
  signal array_obj_ref_1131_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1131_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1131_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1131_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1473_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1131_final_reg_req_0 : boolean;
  signal array_obj_ref_1131_final_reg_ack_0 : boolean;
  signal type_cast_1412_inst_req_0 : boolean;
  signal array_obj_ref_1446_index_0_resize_req_0 : boolean;
  signal binary_1466_inst_req_1 : boolean;
  signal type_cast_1412_inst_ack_0 : boolean;
  signal array_obj_ref_1446_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1446_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1446_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1136_base_resize_req_0 : boolean;
  signal array_obj_ref_1136_base_resize_ack_0 : boolean;
  signal array_obj_ref_1136_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1136_root_address_inst_ack_0 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal array_obj_ref_1136_root_address_inst_req_1 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal array_obj_ref_1136_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1136_final_reg_req_0 : boolean;
  signal array_obj_ref_1136_final_reg_ack_0 : boolean;
  signal array_obj_ref_1446_offset_inst_req_0 : boolean;
  signal array_obj_ref_1446_offset_inst_ack_0 : boolean;
  signal type_cast_1460_inst_req_0 : boolean;
  signal array_obj_ref_1141_base_resize_req_0 : boolean;
  signal array_obj_ref_1141_base_resize_ack_0 : boolean;
  signal array_obj_ref_1470_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1470_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1141_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1141_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1141_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1141_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1141_final_reg_req_0 : boolean;
  signal array_obj_ref_1141_final_reg_ack_0 : boolean;
  signal simple_obj_ref_1152_inst_req_0 : boolean;
  signal simple_obj_ref_1152_inst_ack_0 : boolean;
  signal simple_obj_ref_1161_inst_req_0 : boolean;
  signal simple_obj_ref_1161_inst_ack_0 : boolean;
  signal type_cast_1165_inst_req_0 : boolean;
  signal type_cast_1165_inst_ack_0 : boolean;
  signal switch_stmt_1167_branch_default_req_0 : boolean;
  signal switch_stmt_1167_select_expr_0_req_0 : boolean;
  signal switch_stmt_1167_select_expr_0_ack_0 : boolean;
  signal switch_stmt_1167_select_expr_0_req_1 : boolean;
  signal switch_stmt_1167_select_expr_0_ack_1 : boolean;
  signal switch_stmt_1167_branch_0_req_0 : boolean;
  signal switch_stmt_1167_select_expr_1_req_0 : boolean;
  signal switch_stmt_1167_select_expr_1_ack_0 : boolean;
  signal switch_stmt_1167_select_expr_1_req_1 : boolean;
  signal switch_stmt_1167_select_expr_1_ack_1 : boolean;
  signal switch_stmt_1167_branch_1_req_0 : boolean;
  signal switch_stmt_1167_branch_0_ack_1 : boolean;
  signal switch_stmt_1167_branch_1_ack_1 : boolean;
  signal switch_stmt_1167_branch_default_ack_0 : boolean;
  signal binary_1182_inst_req_0 : boolean;
  signal binary_1182_inst_ack_0 : boolean;
  signal binary_1182_inst_req_1 : boolean;
  signal binary_1182_inst_ack_1 : boolean;
  signal type_cast_1186_inst_req_0 : boolean;
  signal type_cast_1186_inst_ack_0 : boolean;
  signal ptr_deref_1189_base_resize_req_0 : boolean;
  signal ptr_deref_1189_base_resize_ack_0 : boolean;
  signal ptr_deref_1189_root_address_inst_req_0 : boolean;
  signal ptr_deref_1189_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1189_addr_0_req_0 : boolean;
  signal ptr_deref_1189_addr_0_ack_0 : boolean;
  signal ptr_deref_1189_gather_scatter_req_0 : boolean;
  signal ptr_deref_1189_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1189_store_0_req_0 : boolean;
  signal ptr_deref_1189_store_0_ack_0 : boolean;
  signal ptr_deref_1189_store_0_req_1 : boolean;
  signal ptr_deref_1189_store_0_ack_1 : boolean;
  signal binary_1196_inst_req_0 : boolean;
  signal binary_1196_inst_ack_0 : boolean;
  signal binary_1196_inst_req_1 : boolean;
  signal binary_1196_inst_ack_1 : boolean;
  signal type_cast_1200_inst_req_0 : boolean;
  signal type_cast_1200_inst_ack_0 : boolean;
  signal ptr_deref_1203_base_resize_req_0 : boolean;
  signal ptr_deref_1203_base_resize_ack_0 : boolean;
  signal ptr_deref_1203_root_address_inst_req_0 : boolean;
  signal ptr_deref_1203_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1203_addr_0_req_0 : boolean;
  signal ptr_deref_1203_addr_0_ack_0 : boolean;
  signal ptr_deref_1203_gather_scatter_req_0 : boolean;
  signal ptr_deref_1203_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1203_store_0_req_0 : boolean;
  signal ptr_deref_1203_store_0_ack_0 : boolean;
  signal ptr_deref_1203_store_0_req_1 : boolean;
  signal ptr_deref_1203_store_0_ack_1 : boolean;
  signal binary_1210_inst_req_0 : boolean;
  signal binary_1210_inst_ack_0 : boolean;
  signal binary_1210_inst_req_1 : boolean;
  signal binary_1210_inst_ack_1 : boolean;
  signal type_cast_1294_inst_ack_0 : boolean;
  signal ptr_deref_1425_base_resize_ack_0 : boolean;
  signal ptr_deref_1425_base_resize_req_0 : boolean;
  signal ptr_deref_1449_addr_0_ack_0 : boolean;
  signal ptr_deref_1297_base_resize_req_0 : boolean;
  signal ptr_deref_1297_base_resize_ack_0 : boolean;
  signal ptr_deref_1297_root_address_inst_req_0 : boolean;
  signal ptr_deref_1449_addr_0_req_0 : boolean;
  signal ptr_deref_1297_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1297_addr_0_req_0 : boolean;
  signal array_obj_ref_1446_root_address_inst_req_1 : boolean;
  signal ptr_deref_1297_addr_0_ack_0 : boolean;
  signal array_obj_ref_1470_offset_inst_req_0 : boolean;
  signal ptr_deref_1297_gather_scatter_req_0 : boolean;
  signal ptr_deref_1297_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1297_store_0_req_0 : boolean;
  signal ptr_deref_1297_store_0_ack_0 : boolean;
  signal array_obj_ref_1470_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1470_root_address_inst_req_1 : boolean;
  signal ptr_deref_1297_store_0_req_1 : boolean;
  signal ptr_deref_1297_store_0_ack_1 : boolean;
  signal ptr_deref_1473_store_0_ack_0 : boolean;
  signal ptr_deref_1473_addr_0_ack_0 : boolean;
  signal ptr_deref_1473_base_resize_ack_0 : boolean;
  signal ptr_deref_1389_store_0_ack_0 : boolean;
  signal ptr_deref_1389_store_0_req_0 : boolean;
  signal array_obj_ref_1470_root_address_inst_ack_0 : boolean;
  signal binary_1304_inst_req_0 : boolean;
  signal binary_1304_inst_ack_0 : boolean;
  signal array_obj_ref_1422_final_reg_ack_0 : boolean;
  signal binary_1304_inst_req_1 : boolean;
  signal binary_1304_inst_ack_1 : boolean;
  signal ptr_deref_1449_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1422_final_reg_req_0 : boolean;
  signal array_obj_ref_1422_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1449_root_address_inst_req_0 : boolean;
  signal type_cast_1308_inst_req_0 : boolean;
  signal type_cast_1308_inst_ack_0 : boolean;
  signal ptr_deref_1473_base_resize_req_0 : boolean;
  signal binary_1456_inst_ack_1 : boolean;
  signal array_obj_ref_1422_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1422_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1422_root_address_inst_req_0 : boolean;
  signal binary_1456_inst_req_1 : boolean;
  signal ptr_deref_1389_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1422_base_resize_ack_0 : boolean;
  signal array_obj_ref_1422_base_resize_req_0 : boolean;
  signal array_obj_ref_1470_root_address_inst_req_0 : boolean;
  signal ptr_deref_1311_base_resize_req_0 : boolean;
  signal ptr_deref_1311_base_resize_ack_0 : boolean;
  signal ptr_deref_1389_gather_scatter_req_0 : boolean;
  signal ptr_deref_1311_root_address_inst_req_0 : boolean;
  signal ptr_deref_1311_root_address_inst_ack_0 : boolean;
  signal binary_1456_inst_ack_0 : boolean;
  signal ptr_deref_1311_addr_0_req_0 : boolean;
  signal ptr_deref_1311_addr_0_ack_0 : boolean;
  signal binary_1456_inst_req_0 : boolean;
  signal ptr_deref_1449_base_resize_ack_0 : boolean;
  signal ptr_deref_1311_gather_scatter_req_0 : boolean;
  signal ptr_deref_1311_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1449_base_resize_req_0 : boolean;
  signal ptr_deref_1311_store_0_req_0 : boolean;
  signal ptr_deref_1311_store_0_ack_0 : boolean;
  signal ptr_deref_1311_store_0_req_1 : boolean;
  signal array_obj_ref_1422_offset_inst_ack_0 : boolean;
  signal ptr_deref_1311_store_0_ack_1 : boolean;
  signal ptr_deref_1473_store_0_req_0 : boolean;
  signal ptr_deref_1473_root_address_inst_req_0 : boolean;
  signal ptr_deref_1389_addr_0_ack_0 : boolean;
  signal array_obj_ref_1422_offset_inst_req_0 : boolean;
  signal array_obj_ref_1422_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1389_addr_0_req_0 : boolean;
  signal array_obj_ref_1422_index_0_rename_req_0 : boolean;
  signal binary_1318_inst_req_0 : boolean;
  signal binary_1318_inst_ack_0 : boolean;
  signal binary_1318_inst_req_1 : boolean;
  signal binary_1318_inst_ack_1 : boolean;
  signal array_obj_ref_1422_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1446_final_reg_ack_0 : boolean;
  signal array_obj_ref_1422_index_0_resize_req_0 : boolean;
  signal ptr_deref_1389_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1389_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1446_final_reg_req_0 : boolean;
  signal type_cast_1322_inst_req_0 : boolean;
  signal type_cast_1322_inst_ack_0 : boolean;
  signal array_obj_ref_1446_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1325_base_resize_req_0 : boolean;
  signal ptr_deref_1325_base_resize_ack_0 : boolean;
  signal ptr_deref_1325_root_address_inst_req_0 : boolean;
  signal ptr_deref_1325_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1325_addr_0_req_0 : boolean;
  signal ptr_deref_1325_addr_0_ack_0 : boolean;
  signal ptr_deref_1325_gather_scatter_req_0 : boolean;
  signal ptr_deref_1325_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1325_store_0_req_0 : boolean;
  signal ptr_deref_1325_store_0_ack_0 : boolean;
  signal ptr_deref_1325_store_0_req_1 : boolean;
  signal ptr_deref_1325_store_0_ack_1 : boolean;
  signal binary_1332_inst_req_0 : boolean;
  signal binary_1332_inst_ack_0 : boolean;
  signal binary_1332_inst_req_1 : boolean;
  signal binary_1332_inst_ack_1 : boolean;
  signal type_cast_1336_inst_req_0 : boolean;
  signal type_cast_1336_inst_ack_0 : boolean;
  signal ptr_deref_1339_base_resize_req_0 : boolean;
  signal ptr_deref_1339_base_resize_ack_0 : boolean;
  signal ptr_deref_1339_root_address_inst_req_0 : boolean;
  signal ptr_deref_1339_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1339_addr_0_req_0 : boolean;
  signal ptr_deref_1339_addr_0_ack_0 : boolean;
  signal ptr_deref_1339_gather_scatter_req_0 : boolean;
  signal ptr_deref_1339_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1339_store_0_req_0 : boolean;
  signal ptr_deref_1339_store_0_ack_0 : boolean;
  signal ptr_deref_1339_store_0_req_1 : boolean;
  signal ptr_deref_1339_store_0_ack_1 : boolean;
  signal binary_1346_inst_req_0 : boolean;
  signal binary_1346_inst_ack_0 : boolean;
  signal binary_1346_inst_req_1 : boolean;
  signal binary_1346_inst_ack_1 : boolean;
  signal type_cast_1350_inst_req_0 : boolean;
  signal type_cast_1350_inst_ack_0 : boolean;
  signal ptr_deref_1353_base_resize_req_0 : boolean;
  signal ptr_deref_1353_base_resize_ack_0 : boolean;
  signal ptr_deref_1353_root_address_inst_req_0 : boolean;
  signal ptr_deref_1353_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1353_addr_0_req_0 : boolean;
  signal ptr_deref_1353_addr_0_ack_0 : boolean;
  signal ptr_deref_1353_gather_scatter_req_0 : boolean;
  signal ptr_deref_1353_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1353_store_0_req_0 : boolean;
  signal ptr_deref_1353_store_0_ack_0 : boolean;
  signal ptr_deref_1353_store_0_req_1 : boolean;
  signal ptr_deref_1353_store_0_ack_1 : boolean;
  signal binary_1360_inst_req_0 : boolean;
  signal binary_1360_inst_ack_0 : boolean;
  signal binary_1360_inst_req_1 : boolean;
  signal binary_1360_inst_ack_1 : boolean;
  signal type_cast_1364_inst_req_0 : boolean;
  signal type_cast_1364_inst_ack_0 : boolean;
  signal ptr_deref_1367_base_resize_req_0 : boolean;
  signal ptr_deref_1367_base_resize_ack_0 : boolean;
  signal ptr_deref_1367_root_address_inst_req_0 : boolean;
  signal ptr_deref_1367_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1367_addr_0_req_0 : boolean;
  signal ptr_deref_1367_addr_0_ack_0 : boolean;
  signal ptr_deref_1367_gather_scatter_req_0 : boolean;
  signal ptr_deref_1367_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1367_store_0_req_0 : boolean;
  signal ptr_deref_1367_store_0_ack_0 : boolean;
  signal ptr_deref_1367_store_0_req_1 : boolean;
  signal ptr_deref_1367_store_0_ack_1 : boolean;
  signal binary_1374_inst_req_0 : boolean;
  signal binary_1374_inst_ack_0 : boolean;
  signal binary_1374_inst_req_1 : boolean;
  signal binary_1374_inst_ack_1 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal ptr_deref_1473_store_0_req_1 : boolean;
  signal ptr_deref_1473_store_0_ack_1 : boolean;
  signal binary_1480_inst_req_0 : boolean;
  signal binary_1480_inst_ack_0 : boolean;
  signal binary_1480_inst_req_1 : boolean;
  signal binary_1480_inst_ack_1 : boolean;
  signal type_cast_1484_inst_req_0 : boolean;
  signal type_cast_1484_inst_ack_0 : boolean;
  signal binary_1490_inst_req_0 : boolean;
  signal binary_1490_inst_ack_0 : boolean;
  signal binary_1490_inst_req_1 : boolean;
  signal binary_1490_inst_ack_1 : boolean;
  signal array_obj_ref_1494_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1494_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1494_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1494_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1494_offset_inst_req_0 : boolean;
  signal array_obj_ref_1494_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1494_base_resize_req_0 : boolean;
  signal array_obj_ref_1494_base_resize_ack_0 : boolean;
  signal array_obj_ref_1494_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1494_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1494_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1494_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1494_final_reg_req_0 : boolean;
  signal array_obj_ref_1494_final_reg_ack_0 : boolean;
  signal ptr_deref_1497_base_resize_req_0 : boolean;
  signal ptr_deref_1497_base_resize_ack_0 : boolean;
  signal ptr_deref_1497_root_address_inst_req_0 : boolean;
  signal ptr_deref_1497_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1497_addr_0_req_0 : boolean;
  signal ptr_deref_1497_addr_0_ack_0 : boolean;
  signal ptr_deref_1497_gather_scatter_req_0 : boolean;
  signal ptr_deref_1497_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1497_store_0_req_0 : boolean;
  signal ptr_deref_1497_store_0_ack_0 : boolean;
  signal ptr_deref_1497_store_0_req_1 : boolean;
  signal ptr_deref_1497_store_0_ack_1 : boolean;
  signal binary_1504_inst_req_0 : boolean;
  signal binary_1504_inst_ack_0 : boolean;
  signal binary_1504_inst_req_1 : boolean;
  signal binary_1504_inst_ack_1 : boolean;
  signal type_cast_1508_inst_req_0 : boolean;
  signal type_cast_1508_inst_ack_0 : boolean;
  signal binary_1514_inst_req_0 : boolean;
  signal binary_1514_inst_ack_0 : boolean;
  signal binary_1514_inst_req_1 : boolean;
  signal binary_1514_inst_ack_1 : boolean;
  signal array_obj_ref_1518_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1518_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1518_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1518_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1518_offset_inst_req_0 : boolean;
  signal array_obj_ref_1518_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1518_base_resize_req_0 : boolean;
  signal array_obj_ref_1518_base_resize_ack_0 : boolean;
  signal array_obj_ref_1518_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1518_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1518_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1518_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1518_final_reg_req_0 : boolean;
  signal array_obj_ref_1518_final_reg_ack_0 : boolean;
  signal ptr_deref_1521_base_resize_req_0 : boolean;
  signal ptr_deref_1521_base_resize_ack_0 : boolean;
  signal ptr_deref_1521_root_address_inst_req_0 : boolean;
  signal ptr_deref_1521_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1521_addr_0_req_0 : boolean;
  signal ptr_deref_1521_addr_0_ack_0 : boolean;
  signal ptr_deref_1521_gather_scatter_req_0 : boolean;
  signal ptr_deref_1521_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1521_store_0_req_0 : boolean;
  signal ptr_deref_1521_store_0_ack_0 : boolean;
  signal ptr_deref_1521_store_0_req_1 : boolean;
  signal ptr_deref_1521_store_0_ack_1 : boolean;
  signal binary_1528_inst_req_0 : boolean;
  signal binary_1528_inst_ack_0 : boolean;
  signal binary_1528_inst_req_1 : boolean;
  signal binary_1528_inst_ack_1 : boolean;
  signal type_cast_1532_inst_req_0 : boolean;
  signal type_cast_1532_inst_ack_0 : boolean;
  signal binary_1538_inst_req_0 : boolean;
  signal binary_1538_inst_ack_0 : boolean;
  signal binary_1538_inst_req_1 : boolean;
  signal binary_1538_inst_ack_1 : boolean;
  signal array_obj_ref_1542_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1542_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1542_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1542_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1542_offset_inst_req_0 : boolean;
  signal array_obj_ref_1542_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1542_base_resize_req_0 : boolean;
  signal array_obj_ref_1542_base_resize_ack_0 : boolean;
  signal array_obj_ref_1542_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1542_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1542_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1542_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1542_final_reg_req_0 : boolean;
  signal array_obj_ref_1542_final_reg_ack_0 : boolean;
  signal ptr_deref_1545_base_resize_req_0 : boolean;
  signal ptr_deref_1545_base_resize_ack_0 : boolean;
  signal ptr_deref_1545_root_address_inst_req_0 : boolean;
  signal ptr_deref_1545_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1545_addr_0_req_0 : boolean;
  signal ptr_deref_1545_addr_0_ack_0 : boolean;
  signal ptr_deref_1545_gather_scatter_req_0 : boolean;
  signal ptr_deref_1545_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1545_store_0_req_0 : boolean;
  signal ptr_deref_1545_store_0_ack_0 : boolean;
  signal ptr_deref_1545_store_0_req_1 : boolean;
  signal ptr_deref_1545_store_0_ack_1 : boolean;
  signal binary_1552_inst_req_0 : boolean;
  signal binary_1552_inst_ack_0 : boolean;
  signal binary_1552_inst_req_1 : boolean;
  signal binary_1552_inst_ack_1 : boolean;
  signal type_cast_1556_inst_req_0 : boolean;
  signal type_cast_1556_inst_ack_0 : boolean;
  signal binary_1562_inst_req_0 : boolean;
  signal binary_1562_inst_ack_0 : boolean;
  signal binary_1562_inst_req_1 : boolean;
  signal binary_1562_inst_ack_1 : boolean;
  signal array_obj_ref_1566_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1566_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1566_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1566_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1566_offset_inst_req_0 : boolean;
  signal array_obj_ref_1566_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1566_base_resize_req_0 : boolean;
  signal array_obj_ref_1566_base_resize_ack_0 : boolean;
  signal array_obj_ref_1566_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1566_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1566_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1566_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1566_final_reg_req_0 : boolean;
  signal array_obj_ref_1566_final_reg_ack_0 : boolean;
  signal ptr_deref_1569_base_resize_req_0 : boolean;
  signal ptr_deref_1569_base_resize_ack_0 : boolean;
  signal ptr_deref_1569_root_address_inst_req_0 : boolean;
  signal ptr_deref_1569_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1569_addr_0_req_0 : boolean;
  signal ptr_deref_1569_addr_0_ack_0 : boolean;
  signal ptr_deref_1569_gather_scatter_req_0 : boolean;
  signal ptr_deref_1569_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1569_store_0_req_0 : boolean;
  signal ptr_deref_1569_store_0_ack_0 : boolean;
  signal ptr_deref_1569_store_0_req_1 : boolean;
  signal ptr_deref_1569_store_0_ack_1 : boolean;
  signal type_cast_1574_inst_req_0 : boolean;
  signal type_cast_1574_inst_ack_0 : boolean;
  signal binary_1580_inst_req_0 : boolean;
  signal binary_1580_inst_ack_0 : boolean;
  signal binary_1580_inst_req_1 : boolean;
  signal binary_1580_inst_ack_1 : boolean;
  signal array_obj_ref_1584_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1584_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1584_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1584_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1584_offset_inst_req_0 : boolean;
  signal array_obj_ref_1584_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1584_base_resize_req_0 : boolean;
  signal array_obj_ref_1584_base_resize_ack_0 : boolean;
  signal array_obj_ref_1584_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1584_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1584_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1584_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1584_final_reg_req_0 : boolean;
  signal array_obj_ref_1584_final_reg_ack_0 : boolean;
  signal ptr_deref_1587_base_resize_req_0 : boolean;
  signal ptr_deref_1587_base_resize_ack_0 : boolean;
  signal ptr_deref_1587_root_address_inst_req_0 : boolean;
  signal ptr_deref_1587_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1587_addr_0_req_0 : boolean;
  signal ptr_deref_1587_addr_0_ack_0 : boolean;
  signal ptr_deref_1587_gather_scatter_req_0 : boolean;
  signal ptr_deref_1587_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1587_store_0_req_0 : boolean;
  signal ptr_deref_1587_store_0_ack_0 : boolean;
  signal ptr_deref_1587_store_0_req_1 : boolean;
  signal ptr_deref_1587_store_0_ack_1 : boolean;
  signal simple_obj_ref_1596_inst_req_0 : boolean;
  signal simple_obj_ref_1596_inst_ack_0 : boolean;
  signal phi_stmt_1071_req_0 : boolean;
  signal type_cast_1077_inst_req_0 : boolean;
  signal type_cast_1077_inst_ack_0 : boolean;
  signal phi_stmt_1071_req_1 : boolean;
  signal phi_stmt_1071_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_input_CP_4300: Block -- control-path 
    signal cp_elements: BooleanArray(786 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(18);
    cp_elements(3) <= OrReduce(cp_elements(33) & cp_elements(778));
    simple_obj_ref_1014_inst_req_0 <= cp_elements(3);
    cp_elements(4) <= cp_elements(105);
    phi_stmt_1071_req_0 <= cp_elements(4);
    cp_elements(5) <= cp_elements(194);
    cp_elements(6) <= OrReduce(cp_elements(216) & cp_elements(786));
    cp_elements(7) <= cp_elements(361);
    cp_elements(8) <= cp_elements(507);
    type_cast_1077_inst_req_0 <= cp_elements(8);
    cp_elements(9) <= cp_elements(773);
    simple_obj_ref_1596_inst_req_0 <= cp_elements(9);
    cp_elements(10) <= cp_elements(0);
    cp_elements(11) <= cp_elements(10);
    cpelement_group_12 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(14));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(12),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_969_gather_scatter_req_0 <= cp_elements(12);
    cp_elements(13) <= cp_elements(10);
    cp_elements(14) <= cp_elements(10);
    cp_elements(15) <= ptr_deref_969_gather_scatter_ack_0;
    ptr_deref_969_store_0_req_0 <= cp_elements(15);
    cp_elements(16) <= ptr_deref_969_store_0_ack_0;
    ptr_deref_969_store_0_req_1 <= cp_elements(16);
    cp_elements(17) <= ptr_deref_969_store_0_ack_1;
    cpelement_group_18 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(13) & cp_elements(17));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(18),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(19) <= simple_obj_ref_981_inst_ack_0;
    simple_obj_ref_992_inst_req_0 <= cp_elements(19);
    cp_elements(20) <= simple_obj_ref_992_inst_ack_0;
    cp_elements(21) <= cp_elements(20);
    cpelement_group_22 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(23) & cp_elements(24));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(22),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_998_inst_req_0 <= cp_elements(22);
    cp_elements(23) <= cp_elements(21);
    cp_elements(24) <= cp_elements(21);
    cp_elements(25) <= binary_998_inst_ack_0;
    binary_998_inst_req_1 <= cp_elements(25);
    cp_elements(26) <= binary_998_inst_ack_1;
    cp_elements(27) <= cp_elements(26);
    cp_elements(28) <= false;
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= cp_elements(26);
    if_stmt_1000_branch_req_0 <= cp_elements(30);
    cp_elements(31) <= cp_elements(30);
    cp_elements(32) <= cp_elements(31);
    cp_elements(33) <= if_stmt_1000_branch_ack_1;
    cp_elements(34) <= cp_elements(31);
    cp_elements(35) <= if_stmt_1000_branch_ack_0;
    cp_elements(36) <= simple_obj_ref_1014_inst_ack_0;
    cp_elements(37) <= cp_elements(36);
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(39) & cp_elements(40));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1018_inst_req_0 <= cp_elements(38);
    cp_elements(39) <= cp_elements(37);
    cp_elements(40) <= cp_elements(37);
    cp_elements(41) <= type_cast_1018_inst_ack_0;
    cpelement_group_42 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(43) & cp_elements(44));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(42),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1023_inst_req_0 <= cp_elements(42);
    cp_elements(43) <= cp_elements(37);
    cp_elements(44) <= cp_elements(37);
    cp_elements(45) <= type_cast_1023_inst_ack_0;
    cp_elements(46) <= cp_elements(37);
    cpelement_group_47 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(46) & cp_elements(51));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(47),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1028_final_reg_req_0 <= cp_elements(47);
    cp_elements(48) <= cp_elements(41);
    array_obj_ref_1028_base_resize_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_1028_base_resize_ack_0;
    array_obj_ref_1028_root_address_inst_req_0 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_1028_root_address_inst_ack_0;
    array_obj_ref_1028_root_address_inst_req_1 <= cp_elements(50);
    cp_elements(51) <= array_obj_ref_1028_root_address_inst_ack_1;
    cp_elements(52) <= array_obj_ref_1028_final_reg_ack_0;
    cp_elements(53) <= cp_elements(37);
    cpelement_group_54 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(58));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(54),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1033_final_reg_req_0 <= cp_elements(54);
    cp_elements(55) <= cp_elements(45);
    array_obj_ref_1033_base_resize_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_1033_base_resize_ack_0;
    array_obj_ref_1033_root_address_inst_req_0 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_1033_root_address_inst_ack_0;
    array_obj_ref_1033_root_address_inst_req_1 <= cp_elements(57);
    cp_elements(58) <= array_obj_ref_1033_root_address_inst_ack_1;
    cp_elements(59) <= array_obj_ref_1033_final_reg_ack_0;
    cp_elements(60) <= cp_elements(37);
    cpelement_group_61 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(65));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(61),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1038_final_reg_req_0 <= cp_elements(61);
    cp_elements(62) <= cp_elements(45);
    array_obj_ref_1038_base_resize_req_0 <= cp_elements(62);
    cp_elements(63) <= array_obj_ref_1038_base_resize_ack_0;
    array_obj_ref_1038_root_address_inst_req_0 <= cp_elements(63);
    cp_elements(64) <= array_obj_ref_1038_root_address_inst_ack_0;
    array_obj_ref_1038_root_address_inst_req_1 <= cp_elements(64);
    cp_elements(65) <= array_obj_ref_1038_root_address_inst_ack_1;
    cp_elements(66) <= array_obj_ref_1038_final_reg_ack_0;
    cp_elements(67) <= cp_elements(37);
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(67) & cp_elements(72));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1043_final_reg_req_0 <= cp_elements(68);
    cp_elements(69) <= cp_elements(45);
    array_obj_ref_1043_base_resize_req_0 <= cp_elements(69);
    cp_elements(70) <= array_obj_ref_1043_base_resize_ack_0;
    array_obj_ref_1043_root_address_inst_req_0 <= cp_elements(70);
    cp_elements(71) <= array_obj_ref_1043_root_address_inst_ack_0;
    array_obj_ref_1043_root_address_inst_req_1 <= cp_elements(71);
    cp_elements(72) <= array_obj_ref_1043_root_address_inst_ack_1;
    cp_elements(73) <= array_obj_ref_1043_final_reg_ack_0;
    cp_elements(74) <= cp_elements(37);
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(74) & cp_elements(79));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1048_final_reg_req_0 <= cp_elements(75);
    cp_elements(76) <= cp_elements(41);
    array_obj_ref_1048_base_resize_req_0 <= cp_elements(76);
    cp_elements(77) <= array_obj_ref_1048_base_resize_ack_0;
    array_obj_ref_1048_root_address_inst_req_0 <= cp_elements(77);
    cp_elements(78) <= array_obj_ref_1048_root_address_inst_ack_0;
    array_obj_ref_1048_root_address_inst_req_1 <= cp_elements(78);
    cp_elements(79) <= array_obj_ref_1048_root_address_inst_ack_1;
    cp_elements(80) <= array_obj_ref_1048_final_reg_ack_0;
    cpelement_group_81 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(80) & cp_elements(82));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(81),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1052_inst_req_0 <= cp_elements(81);
    cp_elements(82) <= cp_elements(37);
    cp_elements(83) <= type_cast_1052_inst_ack_0;
    cp_elements(84) <= cp_elements(37);
    cpelement_group_85 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(84) & cp_elements(89));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(85),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1057_final_reg_req_0 <= cp_elements(85);
    cp_elements(86) <= cp_elements(45);
    array_obj_ref_1057_base_resize_req_0 <= cp_elements(86);
    cp_elements(87) <= array_obj_ref_1057_base_resize_ack_0;
    array_obj_ref_1057_root_address_inst_req_0 <= cp_elements(87);
    cp_elements(88) <= array_obj_ref_1057_root_address_inst_ack_0;
    array_obj_ref_1057_root_address_inst_req_1 <= cp_elements(88);
    cp_elements(89) <= array_obj_ref_1057_root_address_inst_ack_1;
    cp_elements(90) <= array_obj_ref_1057_final_reg_ack_0;
    cp_elements(91) <= cp_elements(37);
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(91) & cp_elements(96));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1062_final_reg_req_0 <= cp_elements(92);
    cp_elements(93) <= cp_elements(45);
    array_obj_ref_1062_base_resize_req_0 <= cp_elements(93);
    cp_elements(94) <= array_obj_ref_1062_base_resize_ack_0;
    array_obj_ref_1062_root_address_inst_req_0 <= cp_elements(94);
    cp_elements(95) <= array_obj_ref_1062_root_address_inst_ack_0;
    array_obj_ref_1062_root_address_inst_req_1 <= cp_elements(95);
    cp_elements(96) <= array_obj_ref_1062_root_address_inst_ack_1;
    cp_elements(97) <= array_obj_ref_1062_final_reg_ack_0;
    cp_elements(98) <= cp_elements(37);
    cpelement_group_99 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(98) & cp_elements(103));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(99),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1067_final_reg_req_0 <= cp_elements(99);
    cp_elements(100) <= cp_elements(45);
    array_obj_ref_1067_base_resize_req_0 <= cp_elements(100);
    cp_elements(101) <= array_obj_ref_1067_base_resize_ack_0;
    array_obj_ref_1067_root_address_inst_req_0 <= cp_elements(101);
    cp_elements(102) <= array_obj_ref_1067_root_address_inst_ack_0;
    array_obj_ref_1067_root_address_inst_req_1 <= cp_elements(102);
    cp_elements(103) <= array_obj_ref_1067_root_address_inst_ack_1;
    cp_elements(104) <= array_obj_ref_1067_final_reg_ack_0;
    cpelement_group_105 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(52) & cp_elements(59) & cp_elements(66) & cp_elements(73) & cp_elements(83) & cp_elements(90) & cp_elements(97) & cp_elements(104));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(105),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(106) <= cp_elements(782);
    cpelement_group_107 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(108) & cp_elements(109));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(107),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1083_inst_req_0 <= cp_elements(107);
    cp_elements(108) <= cp_elements(106);
    cp_elements(109) <= cp_elements(106);
    cp_elements(110) <= binary_1083_inst_ack_0;
    binary_1083_inst_req_1 <= cp_elements(110);
    cp_elements(111) <= binary_1083_inst_ack_1;
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(114));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1089_inst_req_0 <= cp_elements(112);
    cp_elements(113) <= cp_elements(106);
    cp_elements(114) <= cp_elements(111);
    cp_elements(115) <= binary_1089_inst_ack_0;
    binary_1089_inst_req_1 <= cp_elements(115);
    cp_elements(116) <= binary_1089_inst_ack_1;
    array_obj_ref_1093_index_0_resize_req_0 <= cp_elements(116);
    cp_elements(117) <= cp_elements(106);
    cpelement_group_118 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(117) & cp_elements(127));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1093_final_reg_req_0 <= cp_elements(118);
    cp_elements(119) <= cp_elements(106);
    array_obj_ref_1093_base_resize_req_0 <= cp_elements(119);
    cp_elements(120) <= array_obj_ref_1093_index_0_resize_ack_0;
    array_obj_ref_1093_index_0_scale_req_0 <= cp_elements(120);
    cp_elements(121) <= array_obj_ref_1093_index_0_scale_ack_0;
    array_obj_ref_1093_index_0_scale_req_1 <= cp_elements(121);
    cp_elements(122) <= array_obj_ref_1093_index_0_scale_ack_1;
    array_obj_ref_1093_offset_inst_req_0 <= cp_elements(122);
    cp_elements(123) <= array_obj_ref_1093_offset_inst_ack_0;
    cp_elements(124) <= array_obj_ref_1093_base_resize_ack_0;
    cpelement_group_125 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(123) & cp_elements(124));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(125),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1093_root_address_inst_req_0 <= cp_elements(125);
    cp_elements(126) <= array_obj_ref_1093_root_address_inst_ack_0;
    array_obj_ref_1093_root_address_inst_req_1 <= cp_elements(126);
    cp_elements(127) <= array_obj_ref_1093_root_address_inst_ack_1;
    cp_elements(128) <= array_obj_ref_1093_final_reg_ack_0;
    cpelement_group_129 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(128) & cp_elements(130));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(129),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1097_inst_req_0 <= cp_elements(129);
    cp_elements(130) <= cp_elements(106);
    cp_elements(131) <= type_cast_1097_inst_ack_0;
    cp_elements(132) <= cp_elements(106);
    cpelement_group_133 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(132) & cp_elements(137));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(133),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1102_final_reg_req_0 <= cp_elements(133);
    cp_elements(134) <= cp_elements(131);
    array_obj_ref_1102_base_resize_req_0 <= cp_elements(134);
    cp_elements(135) <= array_obj_ref_1102_base_resize_ack_0;
    array_obj_ref_1102_root_address_inst_req_0 <= cp_elements(135);
    cp_elements(136) <= array_obj_ref_1102_root_address_inst_ack_0;
    array_obj_ref_1102_root_address_inst_req_1 <= cp_elements(136);
    cp_elements(137) <= array_obj_ref_1102_root_address_inst_ack_1;
    cp_elements(138) <= array_obj_ref_1102_final_reg_ack_0;
    cp_elements(139) <= cp_elements(106);
    cpelement_group_140 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(144));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(140),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1107_final_reg_req_0 <= cp_elements(140);
    cp_elements(141) <= cp_elements(131);
    array_obj_ref_1107_base_resize_req_0 <= cp_elements(141);
    cp_elements(142) <= array_obj_ref_1107_base_resize_ack_0;
    array_obj_ref_1107_root_address_inst_req_0 <= cp_elements(142);
    cp_elements(143) <= array_obj_ref_1107_root_address_inst_ack_0;
    array_obj_ref_1107_root_address_inst_req_1 <= cp_elements(143);
    cp_elements(144) <= array_obj_ref_1107_root_address_inst_ack_1;
    cp_elements(145) <= array_obj_ref_1107_final_reg_ack_0;
    cp_elements(146) <= cp_elements(106);
    cpelement_group_147 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(146) & cp_elements(151));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1112_final_reg_req_0 <= cp_elements(147);
    cp_elements(148) <= cp_elements(131);
    array_obj_ref_1112_base_resize_req_0 <= cp_elements(148);
    cp_elements(149) <= array_obj_ref_1112_base_resize_ack_0;
    array_obj_ref_1112_root_address_inst_req_0 <= cp_elements(149);
    cp_elements(150) <= array_obj_ref_1112_root_address_inst_ack_0;
    array_obj_ref_1112_root_address_inst_req_1 <= cp_elements(150);
    cp_elements(151) <= array_obj_ref_1112_root_address_inst_ack_1;
    cp_elements(152) <= array_obj_ref_1112_final_reg_ack_0;
    cpelement_group_153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(154) & cp_elements(155));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1118_inst_req_0 <= cp_elements(153);
    cp_elements(154) <= cp_elements(106);
    cp_elements(155) <= cp_elements(111);
    cp_elements(156) <= binary_1118_inst_ack_0;
    binary_1118_inst_req_1 <= cp_elements(156);
    cp_elements(157) <= binary_1118_inst_ack_1;
    array_obj_ref_1122_index_0_resize_req_0 <= cp_elements(157);
    cp_elements(158) <= cp_elements(106);
    cpelement_group_159 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(158) & cp_elements(168));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(159),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1122_final_reg_req_0 <= cp_elements(159);
    cp_elements(160) <= cp_elements(106);
    array_obj_ref_1122_base_resize_req_0 <= cp_elements(160);
    cp_elements(161) <= array_obj_ref_1122_index_0_resize_ack_0;
    array_obj_ref_1122_index_0_scale_req_0 <= cp_elements(161);
    cp_elements(162) <= array_obj_ref_1122_index_0_scale_ack_0;
    array_obj_ref_1122_index_0_scale_req_1 <= cp_elements(162);
    cp_elements(163) <= array_obj_ref_1122_index_0_scale_ack_1;
    array_obj_ref_1122_offset_inst_req_0 <= cp_elements(163);
    cp_elements(164) <= array_obj_ref_1122_offset_inst_ack_0;
    cp_elements(165) <= array_obj_ref_1122_base_resize_ack_0;
    cpelement_group_166 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(164) & cp_elements(165));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(166),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1122_root_address_inst_req_0 <= cp_elements(166);
    cp_elements(167) <= array_obj_ref_1122_root_address_inst_ack_0;
    array_obj_ref_1122_root_address_inst_req_1 <= cp_elements(167);
    cp_elements(168) <= array_obj_ref_1122_root_address_inst_ack_1;
    cp_elements(169) <= array_obj_ref_1122_final_reg_ack_0;
    cpelement_group_170 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(171));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(170),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1126_inst_req_0 <= cp_elements(170);
    cp_elements(171) <= cp_elements(106);
    cp_elements(172) <= type_cast_1126_inst_ack_0;
    cp_elements(173) <= cp_elements(106);
    cpelement_group_174 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(173) & cp_elements(178));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(174),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1131_final_reg_req_0 <= cp_elements(174);
    cp_elements(175) <= cp_elements(172);
    array_obj_ref_1131_base_resize_req_0 <= cp_elements(175);
    cp_elements(176) <= array_obj_ref_1131_base_resize_ack_0;
    array_obj_ref_1131_root_address_inst_req_0 <= cp_elements(176);
    cp_elements(177) <= array_obj_ref_1131_root_address_inst_ack_0;
    array_obj_ref_1131_root_address_inst_req_1 <= cp_elements(177);
    cp_elements(178) <= array_obj_ref_1131_root_address_inst_ack_1;
    cp_elements(179) <= array_obj_ref_1131_final_reg_ack_0;
    cp_elements(180) <= cp_elements(106);
    cpelement_group_181 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(180) & cp_elements(185));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(181),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1136_final_reg_req_0 <= cp_elements(181);
    cp_elements(182) <= cp_elements(172);
    array_obj_ref_1136_base_resize_req_0 <= cp_elements(182);
    cp_elements(183) <= array_obj_ref_1136_base_resize_ack_0;
    array_obj_ref_1136_root_address_inst_req_0 <= cp_elements(183);
    cp_elements(184) <= array_obj_ref_1136_root_address_inst_ack_0;
    array_obj_ref_1136_root_address_inst_req_1 <= cp_elements(184);
    cp_elements(185) <= array_obj_ref_1136_root_address_inst_ack_1;
    cp_elements(186) <= array_obj_ref_1136_final_reg_ack_0;
    cp_elements(187) <= cp_elements(106);
    cpelement_group_188 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(187) & cp_elements(192));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(188),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1141_final_reg_req_0 <= cp_elements(188);
    cp_elements(189) <= cp_elements(172);
    array_obj_ref_1141_base_resize_req_0 <= cp_elements(189);
    cp_elements(190) <= array_obj_ref_1141_base_resize_ack_0;
    array_obj_ref_1141_root_address_inst_req_0 <= cp_elements(190);
    cp_elements(191) <= array_obj_ref_1141_root_address_inst_ack_0;
    array_obj_ref_1141_root_address_inst_req_1 <= cp_elements(191);
    cp_elements(192) <= array_obj_ref_1141_root_address_inst_ack_1;
    cp_elements(193) <= array_obj_ref_1141_final_reg_ack_0;
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(5 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(138) & cp_elements(145) & cp_elements(152) & cp_elements(179) & cp_elements(186) & cp_elements(193));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(195) <= simple_obj_ref_1152_inst_ack_0;
    simple_obj_ref_1161_inst_req_0 <= cp_elements(195);
    cp_elements(196) <= simple_obj_ref_1161_inst_ack_0;
    cp_elements(197) <= cp_elements(196);
    cpelement_group_198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(199) & cp_elements(200));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1165_inst_req_0 <= cp_elements(198);
    cp_elements(199) <= cp_elements(197);
    cp_elements(200) <= cp_elements(197);
    cp_elements(201) <= type_cast_1165_inst_ack_0;
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= false;
    cp_elements(204) <= cp_elements(203);
    cp_elements(205) <= cp_elements(201);
    cp_elements(206) <= cp_elements(205);
    cp_elements(207) <= cp_elements(206);
    switch_stmt_1167_select_expr_0_req_0 <= cp_elements(207);
    cp_elements(208) <= switch_stmt_1167_select_expr_0_ack_0;
    switch_stmt_1167_select_expr_0_req_1 <= cp_elements(208);
    cp_elements(209) <= switch_stmt_1167_select_expr_0_ack_1;
    switch_stmt_1167_branch_0_req_0 <= cp_elements(209);
    cp_elements(210) <= cp_elements(206);
    switch_stmt_1167_select_expr_1_req_0 <= cp_elements(210);
    cp_elements(211) <= switch_stmt_1167_select_expr_1_ack_0;
    switch_stmt_1167_select_expr_1_req_1 <= cp_elements(211);
    cp_elements(212) <= switch_stmt_1167_select_expr_1_ack_1;
    switch_stmt_1167_branch_1_req_0 <= cp_elements(212);
    cpelement_group_213 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(209) & cp_elements(212));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(213),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    switch_stmt_1167_branch_default_req_0 <= cp_elements(213);
    cp_elements(214) <= cp_elements(213);
    cp_elements(215) <= cp_elements(214);
    cp_elements(216) <= switch_stmt_1167_branch_0_ack_1;
    cp_elements(217) <= cp_elements(214);
    cp_elements(218) <= switch_stmt_1167_branch_1_ack_1;
    cp_elements(219) <= cp_elements(214);
    cp_elements(220) <= switch_stmt_1167_branch_default_ack_0;
    cp_elements(221) <= cp_elements(6);
    cpelement_group_222 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(224));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(222),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1182_inst_req_0 <= cp_elements(222);
    cp_elements(223) <= cp_elements(221);
    cp_elements(224) <= cp_elements(221);
    cp_elements(225) <= binary_1182_inst_ack_0;
    binary_1182_inst_req_1 <= cp_elements(225);
    cp_elements(226) <= binary_1182_inst_ack_1;
    cpelement_group_227 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(226) & cp_elements(228));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(227),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1186_inst_req_0 <= cp_elements(227);
    cp_elements(228) <= cp_elements(221);
    cp_elements(229) <= type_cast_1186_inst_ack_0;
    cpelement_group_230 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(229) & cp_elements(231) & cp_elements(235));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(230),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1189_gather_scatter_req_0 <= cp_elements(230);
    cp_elements(231) <= cp_elements(221);
    cp_elements(232) <= cp_elements(231);
    ptr_deref_1189_base_resize_req_0 <= cp_elements(232);
    cp_elements(233) <= ptr_deref_1189_base_resize_ack_0;
    ptr_deref_1189_root_address_inst_req_0 <= cp_elements(233);
    cp_elements(234) <= ptr_deref_1189_root_address_inst_ack_0;
    ptr_deref_1189_addr_0_req_0 <= cp_elements(234);
    cp_elements(235) <= ptr_deref_1189_addr_0_ack_0;
    cp_elements(236) <= ptr_deref_1189_gather_scatter_ack_0;
    ptr_deref_1189_store_0_req_0 <= cp_elements(236);
    cp_elements(237) <= ptr_deref_1189_store_0_ack_0;
    cp_elements(238) <= cp_elements(237);
    ptr_deref_1189_store_0_req_1 <= cp_elements(238);
    cp_elements(239) <= ptr_deref_1189_store_0_ack_1;
    cpelement_group_240 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(241) & cp_elements(242));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(240),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1196_inst_req_0 <= cp_elements(240);
    cp_elements(241) <= cp_elements(221);
    cp_elements(242) <= cp_elements(221);
    cp_elements(243) <= binary_1196_inst_ack_0;
    binary_1196_inst_req_1 <= cp_elements(243);
    cp_elements(244) <= binary_1196_inst_ack_1;
    cpelement_group_245 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(244) & cp_elements(246));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(245),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1200_inst_req_0 <= cp_elements(245);
    cp_elements(246) <= cp_elements(221);
    cp_elements(247) <= type_cast_1200_inst_ack_0;
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(237) & cp_elements(247) & cp_elements(249) & cp_elements(253));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1203_gather_scatter_req_0 <= cp_elements(248);
    cp_elements(249) <= cp_elements(221);
    cp_elements(250) <= cp_elements(249);
    ptr_deref_1203_base_resize_req_0 <= cp_elements(250);
    cp_elements(251) <= ptr_deref_1203_base_resize_ack_0;
    ptr_deref_1203_root_address_inst_req_0 <= cp_elements(251);
    cp_elements(252) <= ptr_deref_1203_root_address_inst_ack_0;
    ptr_deref_1203_addr_0_req_0 <= cp_elements(252);
    cp_elements(253) <= ptr_deref_1203_addr_0_ack_0;
    cp_elements(254) <= ptr_deref_1203_gather_scatter_ack_0;
    ptr_deref_1203_store_0_req_0 <= cp_elements(254);
    cp_elements(255) <= ptr_deref_1203_store_0_ack_0;
    cp_elements(256) <= cp_elements(255);
    ptr_deref_1203_store_0_req_1 <= cp_elements(256);
    cp_elements(257) <= ptr_deref_1203_store_0_ack_1;
    cpelement_group_258 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(259) & cp_elements(260));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(258),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1210_inst_req_0 <= cp_elements(258);
    cp_elements(259) <= cp_elements(221);
    cp_elements(260) <= cp_elements(221);
    cp_elements(261) <= binary_1210_inst_ack_0;
    binary_1210_inst_req_1 <= cp_elements(261);
    cp_elements(262) <= binary_1210_inst_ack_1;
    cpelement_group_263 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(264));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(263),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1214_inst_req_0 <= cp_elements(263);
    cp_elements(264) <= cp_elements(221);
    cp_elements(265) <= type_cast_1214_inst_ack_0;
    cpelement_group_266 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(255) & cp_elements(265) & cp_elements(267) & cp_elements(271));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(266),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1217_gather_scatter_req_0 <= cp_elements(266);
    cp_elements(267) <= cp_elements(221);
    cp_elements(268) <= cp_elements(267);
    ptr_deref_1217_base_resize_req_0 <= cp_elements(268);
    cp_elements(269) <= ptr_deref_1217_base_resize_ack_0;
    ptr_deref_1217_root_address_inst_req_0 <= cp_elements(269);
    cp_elements(270) <= ptr_deref_1217_root_address_inst_ack_0;
    ptr_deref_1217_addr_0_req_0 <= cp_elements(270);
    cp_elements(271) <= ptr_deref_1217_addr_0_ack_0;
    cp_elements(272) <= ptr_deref_1217_gather_scatter_ack_0;
    ptr_deref_1217_store_0_req_0 <= cp_elements(272);
    cp_elements(273) <= ptr_deref_1217_store_0_ack_0;
    cp_elements(274) <= cp_elements(273);
    ptr_deref_1217_store_0_req_1 <= cp_elements(274);
    cp_elements(275) <= ptr_deref_1217_store_0_ack_1;
    cpelement_group_276 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(277) & cp_elements(278));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(276),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1224_inst_req_0 <= cp_elements(276);
    cp_elements(277) <= cp_elements(221);
    cp_elements(278) <= cp_elements(221);
    cp_elements(279) <= binary_1224_inst_ack_0;
    binary_1224_inst_req_1 <= cp_elements(279);
    cp_elements(280) <= binary_1224_inst_ack_1;
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(280) & cp_elements(282));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1228_inst_req_0 <= cp_elements(281);
    cp_elements(282) <= cp_elements(221);
    cp_elements(283) <= type_cast_1228_inst_ack_0;
    cpelement_group_284 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(273) & cp_elements(283) & cp_elements(285) & cp_elements(289));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(284),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1231_gather_scatter_req_0 <= cp_elements(284);
    cp_elements(285) <= cp_elements(221);
    cp_elements(286) <= cp_elements(285);
    ptr_deref_1231_base_resize_req_0 <= cp_elements(286);
    cp_elements(287) <= ptr_deref_1231_base_resize_ack_0;
    ptr_deref_1231_root_address_inst_req_0 <= cp_elements(287);
    cp_elements(288) <= ptr_deref_1231_root_address_inst_ack_0;
    ptr_deref_1231_addr_0_req_0 <= cp_elements(288);
    cp_elements(289) <= ptr_deref_1231_addr_0_ack_0;
    cp_elements(290) <= ptr_deref_1231_gather_scatter_ack_0;
    ptr_deref_1231_store_0_req_0 <= cp_elements(290);
    cp_elements(291) <= ptr_deref_1231_store_0_ack_0;
    cp_elements(292) <= cp_elements(291);
    ptr_deref_1231_store_0_req_1 <= cp_elements(292);
    cp_elements(293) <= ptr_deref_1231_store_0_ack_1;
    cpelement_group_294 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(295) & cp_elements(296));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(294),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1238_inst_req_0 <= cp_elements(294);
    cp_elements(295) <= cp_elements(221);
    cp_elements(296) <= cp_elements(221);
    cp_elements(297) <= binary_1238_inst_ack_0;
    binary_1238_inst_req_1 <= cp_elements(297);
    cp_elements(298) <= binary_1238_inst_ack_1;
    cpelement_group_299 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(298) & cp_elements(300));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(299),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1242_inst_req_0 <= cp_elements(299);
    cp_elements(300) <= cp_elements(221);
    cp_elements(301) <= type_cast_1242_inst_ack_0;
    cpelement_group_302 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(301) & cp_elements(303) & cp_elements(307));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(302),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1245_gather_scatter_req_0 <= cp_elements(302);
    cp_elements(303) <= cp_elements(221);
    cp_elements(304) <= cp_elements(303);
    ptr_deref_1245_base_resize_req_0 <= cp_elements(304);
    cp_elements(305) <= ptr_deref_1245_base_resize_ack_0;
    ptr_deref_1245_root_address_inst_req_0 <= cp_elements(305);
    cp_elements(306) <= ptr_deref_1245_root_address_inst_ack_0;
    ptr_deref_1245_addr_0_req_0 <= cp_elements(306);
    cp_elements(307) <= ptr_deref_1245_addr_0_ack_0;
    cp_elements(308) <= ptr_deref_1245_gather_scatter_ack_0;
    ptr_deref_1245_store_0_req_0 <= cp_elements(308);
    cp_elements(309) <= ptr_deref_1245_store_0_ack_0;
    cp_elements(310) <= cp_elements(309);
    ptr_deref_1245_store_0_req_1 <= cp_elements(310);
    cp_elements(311) <= ptr_deref_1245_store_0_ack_1;
    cpelement_group_312 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(313) & cp_elements(314));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(312),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1252_inst_req_0 <= cp_elements(312);
    cp_elements(313) <= cp_elements(221);
    cp_elements(314) <= cp_elements(221);
    cp_elements(315) <= binary_1252_inst_ack_0;
    binary_1252_inst_req_1 <= cp_elements(315);
    cp_elements(316) <= binary_1252_inst_ack_1;
    cpelement_group_317 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(316) & cp_elements(318));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(317),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1256_inst_req_0 <= cp_elements(317);
    cp_elements(318) <= cp_elements(221);
    cp_elements(319) <= type_cast_1256_inst_ack_0;
    cpelement_group_320 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(309) & cp_elements(319) & cp_elements(321) & cp_elements(325));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(320),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1259_gather_scatter_req_0 <= cp_elements(320);
    cp_elements(321) <= cp_elements(221);
    cp_elements(322) <= cp_elements(321);
    ptr_deref_1259_base_resize_req_0 <= cp_elements(322);
    cp_elements(323) <= ptr_deref_1259_base_resize_ack_0;
    ptr_deref_1259_root_address_inst_req_0 <= cp_elements(323);
    cp_elements(324) <= ptr_deref_1259_root_address_inst_ack_0;
    ptr_deref_1259_addr_0_req_0 <= cp_elements(324);
    cp_elements(325) <= ptr_deref_1259_addr_0_ack_0;
    cp_elements(326) <= ptr_deref_1259_gather_scatter_ack_0;
    ptr_deref_1259_store_0_req_0 <= cp_elements(326);
    cp_elements(327) <= ptr_deref_1259_store_0_ack_0;
    cp_elements(328) <= cp_elements(327);
    ptr_deref_1259_store_0_req_1 <= cp_elements(328);
    cp_elements(329) <= ptr_deref_1259_store_0_ack_1;
    cpelement_group_330 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(331) & cp_elements(332));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(330),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1266_inst_req_0 <= cp_elements(330);
    cp_elements(331) <= cp_elements(221);
    cp_elements(332) <= cp_elements(221);
    cp_elements(333) <= binary_1266_inst_ack_0;
    binary_1266_inst_req_1 <= cp_elements(333);
    cp_elements(334) <= binary_1266_inst_ack_1;
    cpelement_group_335 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(334) & cp_elements(336));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(335),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1270_inst_req_0 <= cp_elements(335);
    cp_elements(336) <= cp_elements(221);
    cp_elements(337) <= type_cast_1270_inst_ack_0;
    cpelement_group_338 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(327) & cp_elements(337) & cp_elements(339) & cp_elements(343));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(338),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1273_gather_scatter_req_0 <= cp_elements(338);
    cp_elements(339) <= cp_elements(221);
    cp_elements(340) <= cp_elements(339);
    ptr_deref_1273_base_resize_req_0 <= cp_elements(340);
    cp_elements(341) <= ptr_deref_1273_base_resize_ack_0;
    ptr_deref_1273_root_address_inst_req_0 <= cp_elements(341);
    cp_elements(342) <= ptr_deref_1273_root_address_inst_ack_0;
    ptr_deref_1273_addr_0_req_0 <= cp_elements(342);
    cp_elements(343) <= ptr_deref_1273_addr_0_ack_0;
    cp_elements(344) <= ptr_deref_1273_gather_scatter_ack_0;
    ptr_deref_1273_store_0_req_0 <= cp_elements(344);
    cp_elements(345) <= ptr_deref_1273_store_0_ack_0;
    cp_elements(346) <= cp_elements(345);
    ptr_deref_1273_store_0_req_1 <= cp_elements(346);
    cp_elements(347) <= ptr_deref_1273_store_0_ack_1;
    cpelement_group_348 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(349) & cp_elements(350));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(348),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1278_inst_req_0 <= cp_elements(348);
    cp_elements(349) <= cp_elements(221);
    cp_elements(350) <= cp_elements(221);
    cp_elements(351) <= type_cast_1278_inst_ack_0;
    cpelement_group_352 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(345) & cp_elements(351) & cp_elements(353) & cp_elements(357));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(352),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1281_gather_scatter_req_0 <= cp_elements(352);
    cp_elements(353) <= cp_elements(221);
    cp_elements(354) <= cp_elements(353);
    ptr_deref_1281_base_resize_req_0 <= cp_elements(354);
    cp_elements(355) <= ptr_deref_1281_base_resize_ack_0;
    ptr_deref_1281_root_address_inst_req_0 <= cp_elements(355);
    cp_elements(356) <= ptr_deref_1281_root_address_inst_ack_0;
    ptr_deref_1281_addr_0_req_0 <= cp_elements(356);
    cp_elements(357) <= ptr_deref_1281_addr_0_ack_0;
    cp_elements(358) <= ptr_deref_1281_gather_scatter_ack_0;
    ptr_deref_1281_store_0_req_0 <= cp_elements(358);
    cp_elements(359) <= ptr_deref_1281_store_0_ack_0;
    ptr_deref_1281_store_0_req_1 <= cp_elements(359);
    cp_elements(360) <= ptr_deref_1281_store_0_ack_1;
    cpelement_group_361 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(239) & cp_elements(257) & cp_elements(275) & cp_elements(293) & cp_elements(311) & cp_elements(329) & cp_elements(347) & cp_elements(360));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(361),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(362) <= cp_elements(218);
    cpelement_group_363 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(364) & cp_elements(365));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(363),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1290_inst_req_0 <= cp_elements(363);
    cp_elements(364) <= cp_elements(362);
    cp_elements(365) <= cp_elements(362);
    cp_elements(366) <= binary_1290_inst_ack_0;
    binary_1290_inst_req_1 <= cp_elements(366);
    cp_elements(367) <= binary_1290_inst_ack_1;
    cpelement_group_368 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(367) & cp_elements(369));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(368),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1294_inst_req_0 <= cp_elements(368);
    cp_elements(369) <= cp_elements(362);
    cp_elements(370) <= type_cast_1294_inst_ack_0;
    cpelement_group_371 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(370) & cp_elements(372) & cp_elements(376));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(371),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1297_gather_scatter_req_0 <= cp_elements(371);
    cp_elements(372) <= cp_elements(362);
    cp_elements(373) <= cp_elements(372);
    ptr_deref_1297_base_resize_req_0 <= cp_elements(373);
    cp_elements(374) <= ptr_deref_1297_base_resize_ack_0;
    ptr_deref_1297_root_address_inst_req_0 <= cp_elements(374);
    cp_elements(375) <= ptr_deref_1297_root_address_inst_ack_0;
    ptr_deref_1297_addr_0_req_0 <= cp_elements(375);
    cp_elements(376) <= ptr_deref_1297_addr_0_ack_0;
    cp_elements(377) <= ptr_deref_1297_gather_scatter_ack_0;
    ptr_deref_1297_store_0_req_0 <= cp_elements(377);
    cp_elements(378) <= ptr_deref_1297_store_0_ack_0;
    cp_elements(379) <= cp_elements(378);
    ptr_deref_1297_store_0_req_1 <= cp_elements(379);
    cp_elements(380) <= ptr_deref_1297_store_0_ack_1;
    cpelement_group_381 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(382) & cp_elements(383));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(381),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1304_inst_req_0 <= cp_elements(381);
    cp_elements(382) <= cp_elements(362);
    cp_elements(383) <= cp_elements(362);
    cp_elements(384) <= binary_1304_inst_ack_0;
    binary_1304_inst_req_1 <= cp_elements(384);
    cp_elements(385) <= binary_1304_inst_ack_1;
    cpelement_group_386 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(385) & cp_elements(387));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(386),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1308_inst_req_0 <= cp_elements(386);
    cp_elements(387) <= cp_elements(362);
    cp_elements(388) <= type_cast_1308_inst_ack_0;
    cpelement_group_389 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(378) & cp_elements(388) & cp_elements(390) & cp_elements(394));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(389),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1311_gather_scatter_req_0 <= cp_elements(389);
    cp_elements(390) <= cp_elements(362);
    cp_elements(391) <= cp_elements(390);
    ptr_deref_1311_base_resize_req_0 <= cp_elements(391);
    cp_elements(392) <= ptr_deref_1311_base_resize_ack_0;
    ptr_deref_1311_root_address_inst_req_0 <= cp_elements(392);
    cp_elements(393) <= ptr_deref_1311_root_address_inst_ack_0;
    ptr_deref_1311_addr_0_req_0 <= cp_elements(393);
    cp_elements(394) <= ptr_deref_1311_addr_0_ack_0;
    cp_elements(395) <= ptr_deref_1311_gather_scatter_ack_0;
    ptr_deref_1311_store_0_req_0 <= cp_elements(395);
    cp_elements(396) <= ptr_deref_1311_store_0_ack_0;
    cp_elements(397) <= cp_elements(396);
    ptr_deref_1311_store_0_req_1 <= cp_elements(397);
    cp_elements(398) <= ptr_deref_1311_store_0_ack_1;
    cpelement_group_399 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(400) & cp_elements(401));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(399),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1318_inst_req_0 <= cp_elements(399);
    cp_elements(400) <= cp_elements(362);
    cp_elements(401) <= cp_elements(362);
    cp_elements(402) <= binary_1318_inst_ack_0;
    binary_1318_inst_req_1 <= cp_elements(402);
    cp_elements(403) <= binary_1318_inst_ack_1;
    cpelement_group_404 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(403) & cp_elements(405));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(404),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1322_inst_req_0 <= cp_elements(404);
    cp_elements(405) <= cp_elements(362);
    cp_elements(406) <= type_cast_1322_inst_ack_0;
    cpelement_group_407 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(396) & cp_elements(406) & cp_elements(408) & cp_elements(412));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(407),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1325_gather_scatter_req_0 <= cp_elements(407);
    cp_elements(408) <= cp_elements(362);
    cp_elements(409) <= cp_elements(408);
    ptr_deref_1325_base_resize_req_0 <= cp_elements(409);
    cp_elements(410) <= ptr_deref_1325_base_resize_ack_0;
    ptr_deref_1325_root_address_inst_req_0 <= cp_elements(410);
    cp_elements(411) <= ptr_deref_1325_root_address_inst_ack_0;
    ptr_deref_1325_addr_0_req_0 <= cp_elements(411);
    cp_elements(412) <= ptr_deref_1325_addr_0_ack_0;
    cp_elements(413) <= ptr_deref_1325_gather_scatter_ack_0;
    ptr_deref_1325_store_0_req_0 <= cp_elements(413);
    cp_elements(414) <= ptr_deref_1325_store_0_ack_0;
    cp_elements(415) <= cp_elements(414);
    ptr_deref_1325_store_0_req_1 <= cp_elements(415);
    cp_elements(416) <= ptr_deref_1325_store_0_ack_1;
    cpelement_group_417 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(418) & cp_elements(419));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(417),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1332_inst_req_0 <= cp_elements(417);
    cp_elements(418) <= cp_elements(362);
    cp_elements(419) <= cp_elements(362);
    cp_elements(420) <= binary_1332_inst_ack_0;
    binary_1332_inst_req_1 <= cp_elements(420);
    cp_elements(421) <= binary_1332_inst_ack_1;
    cpelement_group_422 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(421) & cp_elements(423));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(422),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1336_inst_req_0 <= cp_elements(422);
    cp_elements(423) <= cp_elements(362);
    cp_elements(424) <= type_cast_1336_inst_ack_0;
    cpelement_group_425 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(414) & cp_elements(424) & cp_elements(426) & cp_elements(430));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(425),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1339_gather_scatter_req_0 <= cp_elements(425);
    cp_elements(426) <= cp_elements(362);
    cp_elements(427) <= cp_elements(426);
    ptr_deref_1339_base_resize_req_0 <= cp_elements(427);
    cp_elements(428) <= ptr_deref_1339_base_resize_ack_0;
    ptr_deref_1339_root_address_inst_req_0 <= cp_elements(428);
    cp_elements(429) <= ptr_deref_1339_root_address_inst_ack_0;
    ptr_deref_1339_addr_0_req_0 <= cp_elements(429);
    cp_elements(430) <= ptr_deref_1339_addr_0_ack_0;
    cp_elements(431) <= ptr_deref_1339_gather_scatter_ack_0;
    ptr_deref_1339_store_0_req_0 <= cp_elements(431);
    cp_elements(432) <= ptr_deref_1339_store_0_ack_0;
    cp_elements(433) <= cp_elements(432);
    ptr_deref_1339_store_0_req_1 <= cp_elements(433);
    cp_elements(434) <= ptr_deref_1339_store_0_ack_1;
    cpelement_group_435 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(436) & cp_elements(437));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(435),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1346_inst_req_0 <= cp_elements(435);
    cp_elements(436) <= cp_elements(362);
    cp_elements(437) <= cp_elements(362);
    cp_elements(438) <= binary_1346_inst_ack_0;
    binary_1346_inst_req_1 <= cp_elements(438);
    cp_elements(439) <= binary_1346_inst_ack_1;
    cpelement_group_440 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(439) & cp_elements(441));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(440),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1350_inst_req_0 <= cp_elements(440);
    cp_elements(441) <= cp_elements(362);
    cp_elements(442) <= type_cast_1350_inst_ack_0;
    cpelement_group_443 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(432) & cp_elements(442) & cp_elements(444) & cp_elements(448));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(443),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1353_gather_scatter_req_0 <= cp_elements(443);
    cp_elements(444) <= cp_elements(362);
    cp_elements(445) <= cp_elements(444);
    ptr_deref_1353_base_resize_req_0 <= cp_elements(445);
    cp_elements(446) <= ptr_deref_1353_base_resize_ack_0;
    ptr_deref_1353_root_address_inst_req_0 <= cp_elements(446);
    cp_elements(447) <= ptr_deref_1353_root_address_inst_ack_0;
    ptr_deref_1353_addr_0_req_0 <= cp_elements(447);
    cp_elements(448) <= ptr_deref_1353_addr_0_ack_0;
    cp_elements(449) <= ptr_deref_1353_gather_scatter_ack_0;
    ptr_deref_1353_store_0_req_0 <= cp_elements(449);
    cp_elements(450) <= ptr_deref_1353_store_0_ack_0;
    cp_elements(451) <= cp_elements(450);
    ptr_deref_1353_store_0_req_1 <= cp_elements(451);
    cp_elements(452) <= ptr_deref_1353_store_0_ack_1;
    cpelement_group_453 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(454) & cp_elements(455));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(453),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1360_inst_req_0 <= cp_elements(453);
    cp_elements(454) <= cp_elements(362);
    cp_elements(455) <= cp_elements(362);
    cp_elements(456) <= binary_1360_inst_ack_0;
    binary_1360_inst_req_1 <= cp_elements(456);
    cp_elements(457) <= binary_1360_inst_ack_1;
    cpelement_group_458 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(457) & cp_elements(459));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(458),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1364_inst_req_0 <= cp_elements(458);
    cp_elements(459) <= cp_elements(362);
    cp_elements(460) <= type_cast_1364_inst_ack_0;
    cpelement_group_461 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(450) & cp_elements(460) & cp_elements(462) & cp_elements(466));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(461),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1367_gather_scatter_req_0 <= cp_elements(461);
    cp_elements(462) <= cp_elements(362);
    cp_elements(463) <= cp_elements(462);
    ptr_deref_1367_base_resize_req_0 <= cp_elements(463);
    cp_elements(464) <= ptr_deref_1367_base_resize_ack_0;
    ptr_deref_1367_root_address_inst_req_0 <= cp_elements(464);
    cp_elements(465) <= ptr_deref_1367_root_address_inst_ack_0;
    ptr_deref_1367_addr_0_req_0 <= cp_elements(465);
    cp_elements(466) <= ptr_deref_1367_addr_0_ack_0;
    cp_elements(467) <= ptr_deref_1367_gather_scatter_ack_0;
    ptr_deref_1367_store_0_req_0 <= cp_elements(467);
    cp_elements(468) <= ptr_deref_1367_store_0_ack_0;
    cp_elements(469) <= cp_elements(468);
    ptr_deref_1367_store_0_req_1 <= cp_elements(469);
    cp_elements(470) <= ptr_deref_1367_store_0_ack_1;
    cpelement_group_471 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(472) & cp_elements(473));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(471),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1374_inst_req_0 <= cp_elements(471);
    cp_elements(472) <= cp_elements(362);
    cp_elements(473) <= cp_elements(362);
    cp_elements(474) <= binary_1374_inst_ack_0;
    binary_1374_inst_req_1 <= cp_elements(474);
    cp_elements(475) <= binary_1374_inst_ack_1;
    cpelement_group_476 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(475) & cp_elements(477));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(476),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1378_inst_req_0 <= cp_elements(476);
    cp_elements(477) <= cp_elements(362);
    cp_elements(478) <= type_cast_1378_inst_ack_0;
    cpelement_group_479 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(468) & cp_elements(478) & cp_elements(480) & cp_elements(484));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(479),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1381_gather_scatter_req_0 <= cp_elements(479);
    cp_elements(480) <= cp_elements(362);
    cp_elements(481) <= cp_elements(480);
    ptr_deref_1381_base_resize_req_0 <= cp_elements(481);
    cp_elements(482) <= ptr_deref_1381_base_resize_ack_0;
    ptr_deref_1381_root_address_inst_req_0 <= cp_elements(482);
    cp_elements(483) <= ptr_deref_1381_root_address_inst_ack_0;
    ptr_deref_1381_addr_0_req_0 <= cp_elements(483);
    cp_elements(484) <= ptr_deref_1381_addr_0_ack_0;
    cp_elements(485) <= ptr_deref_1381_gather_scatter_ack_0;
    ptr_deref_1381_store_0_req_0 <= cp_elements(485);
    cp_elements(486) <= ptr_deref_1381_store_0_ack_0;
    cp_elements(487) <= cp_elements(486);
    ptr_deref_1381_store_0_req_1 <= cp_elements(487);
    cp_elements(488) <= ptr_deref_1381_store_0_ack_1;
    cpelement_group_489 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(490) & cp_elements(491));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(489),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1386_inst_req_0 <= cp_elements(489);
    cp_elements(490) <= cp_elements(362);
    cp_elements(491) <= cp_elements(362);
    cp_elements(492) <= type_cast_1386_inst_ack_0;
    cpelement_group_493 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(486) & cp_elements(492) & cp_elements(494) & cp_elements(498));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(493),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1389_gather_scatter_req_0 <= cp_elements(493);
    cp_elements(494) <= cp_elements(362);
    cp_elements(495) <= cp_elements(494);
    ptr_deref_1389_base_resize_req_0 <= cp_elements(495);
    cp_elements(496) <= ptr_deref_1389_base_resize_ack_0;
    ptr_deref_1389_root_address_inst_req_0 <= cp_elements(496);
    cp_elements(497) <= ptr_deref_1389_root_address_inst_ack_0;
    ptr_deref_1389_addr_0_req_0 <= cp_elements(497);
    cp_elements(498) <= ptr_deref_1389_addr_0_ack_0;
    cp_elements(499) <= ptr_deref_1389_gather_scatter_ack_0;
    ptr_deref_1389_store_0_req_0 <= cp_elements(499);
    cp_elements(500) <= ptr_deref_1389_store_0_ack_0;
    ptr_deref_1389_store_0_req_1 <= cp_elements(500);
    cp_elements(501) <= ptr_deref_1389_store_0_ack_1;
    cpelement_group_502 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(503) & cp_elements(504));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(502),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1396_inst_req_0 <= cp_elements(502);
    cp_elements(503) <= cp_elements(362);
    cp_elements(504) <= cp_elements(362);
    cp_elements(505) <= binary_1396_inst_ack_0;
    binary_1396_inst_req_1 <= cp_elements(505);
    cp_elements(506) <= binary_1396_inst_ack_1;
    cpelement_group_507 : Block -- 
      signal predecessors: BooleanArray(8 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(380) & cp_elements(398) & cp_elements(416) & cp_elements(434) & cp_elements(452) & cp_elements(470) & cp_elements(488) & cp_elements(501) & cp_elements(506));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(507),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(508) <= cp_elements(220);
    cpelement_group_509 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(510) & cp_elements(511));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(509),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1402_inst_req_0 <= cp_elements(509);
    cp_elements(510) <= cp_elements(508);
    cp_elements(511) <= cp_elements(508);
    cp_elements(512) <= type_cast_1402_inst_ack_0;
    cpelement_group_513 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(514) & cp_elements(515));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(513),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1408_inst_req_0 <= cp_elements(513);
    cp_elements(514) <= cp_elements(508);
    cp_elements(515) <= cp_elements(508);
    cp_elements(516) <= binary_1408_inst_ack_0;
    binary_1408_inst_req_1 <= cp_elements(516);
    cp_elements(517) <= binary_1408_inst_ack_1;
    cpelement_group_518 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(517) & cp_elements(519));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(518),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1412_inst_req_0 <= cp_elements(518);
    cp_elements(519) <= cp_elements(508);
    cp_elements(520) <= type_cast_1412_inst_ack_0;
    cpelement_group_521 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(522) & cp_elements(523));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(521),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1418_inst_req_0 <= cp_elements(521);
    cp_elements(522) <= cp_elements(508);
    cp_elements(523) <= cp_elements(508);
    cp_elements(524) <= binary_1418_inst_ack_0;
    binary_1418_inst_req_1 <= cp_elements(524);
    cp_elements(525) <= binary_1418_inst_ack_1;
    cp_elements(526) <= cp_elements(508);
    cpelement_group_527 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(526) & cp_elements(536));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(527),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1422_final_reg_req_0 <= cp_elements(527);
    cp_elements(528) <= cp_elements(512);
    array_obj_ref_1422_base_resize_req_0 <= cp_elements(528);
    cp_elements(529) <= cp_elements(525);
    array_obj_ref_1422_index_0_resize_req_0 <= cp_elements(529);
    cp_elements(530) <= array_obj_ref_1422_index_0_resize_ack_0;
    array_obj_ref_1422_index_0_rename_req_0 <= cp_elements(530);
    cp_elements(531) <= array_obj_ref_1422_index_0_rename_ack_0;
    array_obj_ref_1422_offset_inst_req_0 <= cp_elements(531);
    cp_elements(532) <= array_obj_ref_1422_offset_inst_ack_0;
    cp_elements(533) <= array_obj_ref_1422_base_resize_ack_0;
    cpelement_group_534 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(532) & cp_elements(533));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(534),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1422_root_address_inst_req_0 <= cp_elements(534);
    cp_elements(535) <= array_obj_ref_1422_root_address_inst_ack_0;
    array_obj_ref_1422_root_address_inst_req_1 <= cp_elements(535);
    cp_elements(536) <= array_obj_ref_1422_root_address_inst_ack_1;
    cp_elements(537) <= array_obj_ref_1422_final_reg_ack_0;
    cpelement_group_538 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(520) & cp_elements(537) & cp_elements(542));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(538),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1425_gather_scatter_req_0 <= cp_elements(538);
    cp_elements(539) <= cp_elements(537);
    ptr_deref_1425_base_resize_req_0 <= cp_elements(539);
    cp_elements(540) <= ptr_deref_1425_base_resize_ack_0;
    ptr_deref_1425_root_address_inst_req_0 <= cp_elements(540);
    cp_elements(541) <= ptr_deref_1425_root_address_inst_ack_0;
    ptr_deref_1425_addr_0_req_0 <= cp_elements(541);
    cp_elements(542) <= ptr_deref_1425_addr_0_ack_0;
    cp_elements(543) <= ptr_deref_1425_gather_scatter_ack_0;
    ptr_deref_1425_store_0_req_0 <= cp_elements(543);
    cp_elements(544) <= ptr_deref_1425_store_0_ack_0;
    cp_elements(545) <= cp_elements(544);
    ptr_deref_1425_store_0_req_1 <= cp_elements(545);
    cp_elements(546) <= ptr_deref_1425_store_0_ack_1;
    cpelement_group_547 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(548) & cp_elements(549));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(547),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1432_inst_req_0 <= cp_elements(547);
    cp_elements(548) <= cp_elements(508);
    cp_elements(549) <= cp_elements(508);
    cp_elements(550) <= binary_1432_inst_ack_0;
    binary_1432_inst_req_1 <= cp_elements(550);
    cp_elements(551) <= binary_1432_inst_ack_1;
    cpelement_group_552 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(551) & cp_elements(553));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(552),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1436_inst_req_0 <= cp_elements(552);
    cp_elements(553) <= cp_elements(508);
    cp_elements(554) <= type_cast_1436_inst_ack_0;
    cpelement_group_555 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(556) & cp_elements(557));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(555),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1442_inst_req_0 <= cp_elements(555);
    cp_elements(556) <= cp_elements(508);
    cp_elements(557) <= cp_elements(525);
    cp_elements(558) <= binary_1442_inst_ack_0;
    binary_1442_inst_req_1 <= cp_elements(558);
    cp_elements(559) <= binary_1442_inst_ack_1;
    array_obj_ref_1446_index_0_resize_req_0 <= cp_elements(559);
    cp_elements(560) <= cp_elements(508);
    cpelement_group_561 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(560) & cp_elements(569));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(561),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1446_final_reg_req_0 <= cp_elements(561);
    cp_elements(562) <= cp_elements(512);
    array_obj_ref_1446_base_resize_req_0 <= cp_elements(562);
    cp_elements(563) <= array_obj_ref_1446_index_0_resize_ack_0;
    array_obj_ref_1446_index_0_rename_req_0 <= cp_elements(563);
    cp_elements(564) <= array_obj_ref_1446_index_0_rename_ack_0;
    array_obj_ref_1446_offset_inst_req_0 <= cp_elements(564);
    cp_elements(565) <= array_obj_ref_1446_offset_inst_ack_0;
    cp_elements(566) <= array_obj_ref_1446_base_resize_ack_0;
    cpelement_group_567 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(565) & cp_elements(566));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(567),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1446_root_address_inst_req_0 <= cp_elements(567);
    cp_elements(568) <= array_obj_ref_1446_root_address_inst_ack_0;
    array_obj_ref_1446_root_address_inst_req_1 <= cp_elements(568);
    cp_elements(569) <= array_obj_ref_1446_root_address_inst_ack_1;
    cp_elements(570) <= array_obj_ref_1446_final_reg_ack_0;
    cpelement_group_571 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(544) & cp_elements(554) & cp_elements(570) & cp_elements(575));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(571),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1449_gather_scatter_req_0 <= cp_elements(571);
    cp_elements(572) <= cp_elements(570);
    ptr_deref_1449_base_resize_req_0 <= cp_elements(572);
    cp_elements(573) <= ptr_deref_1449_base_resize_ack_0;
    ptr_deref_1449_root_address_inst_req_0 <= cp_elements(573);
    cp_elements(574) <= ptr_deref_1449_root_address_inst_ack_0;
    ptr_deref_1449_addr_0_req_0 <= cp_elements(574);
    cp_elements(575) <= ptr_deref_1449_addr_0_ack_0;
    cp_elements(576) <= ptr_deref_1449_gather_scatter_ack_0;
    ptr_deref_1449_store_0_req_0 <= cp_elements(576);
    cp_elements(577) <= ptr_deref_1449_store_0_ack_0;
    cp_elements(578) <= cp_elements(577);
    ptr_deref_1449_store_0_req_1 <= cp_elements(578);
    cp_elements(579) <= ptr_deref_1449_store_0_ack_1;
    cpelement_group_580 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(581) & cp_elements(582));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(580),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1456_inst_req_0 <= cp_elements(580);
    cp_elements(581) <= cp_elements(508);
    cp_elements(582) <= cp_elements(508);
    cp_elements(583) <= binary_1456_inst_ack_0;
    binary_1456_inst_req_1 <= cp_elements(583);
    cp_elements(584) <= binary_1456_inst_ack_1;
    cpelement_group_585 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(584) & cp_elements(586));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(585),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1460_inst_req_0 <= cp_elements(585);
    cp_elements(586) <= cp_elements(508);
    cp_elements(587) <= type_cast_1460_inst_ack_0;
    cpelement_group_588 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(589) & cp_elements(590));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(588),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1466_inst_req_0 <= cp_elements(588);
    cp_elements(589) <= cp_elements(508);
    cp_elements(590) <= cp_elements(525);
    cp_elements(591) <= binary_1466_inst_ack_0;
    binary_1466_inst_req_1 <= cp_elements(591);
    cp_elements(592) <= binary_1466_inst_ack_1;
    array_obj_ref_1470_index_0_resize_req_0 <= cp_elements(592);
    cp_elements(593) <= cp_elements(508);
    cpelement_group_594 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(593) & cp_elements(602));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(594),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1470_final_reg_req_0 <= cp_elements(594);
    cp_elements(595) <= cp_elements(512);
    array_obj_ref_1470_base_resize_req_0 <= cp_elements(595);
    cp_elements(596) <= array_obj_ref_1470_index_0_resize_ack_0;
    array_obj_ref_1470_index_0_rename_req_0 <= cp_elements(596);
    cp_elements(597) <= array_obj_ref_1470_index_0_rename_ack_0;
    array_obj_ref_1470_offset_inst_req_0 <= cp_elements(597);
    cp_elements(598) <= array_obj_ref_1470_offset_inst_ack_0;
    cp_elements(599) <= array_obj_ref_1470_base_resize_ack_0;
    cpelement_group_600 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(598) & cp_elements(599));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(600),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1470_root_address_inst_req_0 <= cp_elements(600);
    cp_elements(601) <= array_obj_ref_1470_root_address_inst_ack_0;
    array_obj_ref_1470_root_address_inst_req_1 <= cp_elements(601);
    cp_elements(602) <= array_obj_ref_1470_root_address_inst_ack_1;
    cp_elements(603) <= array_obj_ref_1470_final_reg_ack_0;
    cpelement_group_604 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(577) & cp_elements(587) & cp_elements(603) & cp_elements(608));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(604),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1473_gather_scatter_req_0 <= cp_elements(604);
    cp_elements(605) <= cp_elements(603);
    ptr_deref_1473_base_resize_req_0 <= cp_elements(605);
    cp_elements(606) <= ptr_deref_1473_base_resize_ack_0;
    ptr_deref_1473_root_address_inst_req_0 <= cp_elements(606);
    cp_elements(607) <= ptr_deref_1473_root_address_inst_ack_0;
    ptr_deref_1473_addr_0_req_0 <= cp_elements(607);
    cp_elements(608) <= ptr_deref_1473_addr_0_ack_0;
    cp_elements(609) <= ptr_deref_1473_gather_scatter_ack_0;
    ptr_deref_1473_store_0_req_0 <= cp_elements(609);
    cp_elements(610) <= ptr_deref_1473_store_0_ack_0;
    cp_elements(611) <= cp_elements(610);
    ptr_deref_1473_store_0_req_1 <= cp_elements(611);
    cp_elements(612) <= ptr_deref_1473_store_0_ack_1;
    cpelement_group_613 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(614) & cp_elements(615));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(613),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1480_inst_req_0 <= cp_elements(613);
    cp_elements(614) <= cp_elements(508);
    cp_elements(615) <= cp_elements(508);
    cp_elements(616) <= binary_1480_inst_ack_0;
    binary_1480_inst_req_1 <= cp_elements(616);
    cp_elements(617) <= binary_1480_inst_ack_1;
    cpelement_group_618 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(617) & cp_elements(619));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(618),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1484_inst_req_0 <= cp_elements(618);
    cp_elements(619) <= cp_elements(508);
    cp_elements(620) <= type_cast_1484_inst_ack_0;
    cpelement_group_621 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(622) & cp_elements(623));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(621),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1490_inst_req_0 <= cp_elements(621);
    cp_elements(622) <= cp_elements(508);
    cp_elements(623) <= cp_elements(525);
    cp_elements(624) <= binary_1490_inst_ack_0;
    binary_1490_inst_req_1 <= cp_elements(624);
    cp_elements(625) <= binary_1490_inst_ack_1;
    array_obj_ref_1494_index_0_resize_req_0 <= cp_elements(625);
    cp_elements(626) <= cp_elements(508);
    cpelement_group_627 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(626) & cp_elements(635));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(627),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1494_final_reg_req_0 <= cp_elements(627);
    cp_elements(628) <= cp_elements(512);
    array_obj_ref_1494_base_resize_req_0 <= cp_elements(628);
    cp_elements(629) <= array_obj_ref_1494_index_0_resize_ack_0;
    array_obj_ref_1494_index_0_rename_req_0 <= cp_elements(629);
    cp_elements(630) <= array_obj_ref_1494_index_0_rename_ack_0;
    array_obj_ref_1494_offset_inst_req_0 <= cp_elements(630);
    cp_elements(631) <= array_obj_ref_1494_offset_inst_ack_0;
    cp_elements(632) <= array_obj_ref_1494_base_resize_ack_0;
    cpelement_group_633 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(631) & cp_elements(632));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(633),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1494_root_address_inst_req_0 <= cp_elements(633);
    cp_elements(634) <= array_obj_ref_1494_root_address_inst_ack_0;
    array_obj_ref_1494_root_address_inst_req_1 <= cp_elements(634);
    cp_elements(635) <= array_obj_ref_1494_root_address_inst_ack_1;
    cp_elements(636) <= array_obj_ref_1494_final_reg_ack_0;
    cpelement_group_637 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(610) & cp_elements(620) & cp_elements(636) & cp_elements(641));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(637),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1497_gather_scatter_req_0 <= cp_elements(637);
    cp_elements(638) <= cp_elements(636);
    ptr_deref_1497_base_resize_req_0 <= cp_elements(638);
    cp_elements(639) <= ptr_deref_1497_base_resize_ack_0;
    ptr_deref_1497_root_address_inst_req_0 <= cp_elements(639);
    cp_elements(640) <= ptr_deref_1497_root_address_inst_ack_0;
    ptr_deref_1497_addr_0_req_0 <= cp_elements(640);
    cp_elements(641) <= ptr_deref_1497_addr_0_ack_0;
    cp_elements(642) <= ptr_deref_1497_gather_scatter_ack_0;
    ptr_deref_1497_store_0_req_0 <= cp_elements(642);
    cp_elements(643) <= ptr_deref_1497_store_0_ack_0;
    cp_elements(644) <= cp_elements(643);
    ptr_deref_1497_store_0_req_1 <= cp_elements(644);
    cp_elements(645) <= ptr_deref_1497_store_0_ack_1;
    cpelement_group_646 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(647) & cp_elements(648));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(646),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1504_inst_req_0 <= cp_elements(646);
    cp_elements(647) <= cp_elements(508);
    cp_elements(648) <= cp_elements(508);
    cp_elements(649) <= binary_1504_inst_ack_0;
    binary_1504_inst_req_1 <= cp_elements(649);
    cp_elements(650) <= binary_1504_inst_ack_1;
    cpelement_group_651 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(650) & cp_elements(652));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(651),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1508_inst_req_0 <= cp_elements(651);
    cp_elements(652) <= cp_elements(508);
    cp_elements(653) <= type_cast_1508_inst_ack_0;
    cpelement_group_654 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(655) & cp_elements(656));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(654),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1514_inst_req_0 <= cp_elements(654);
    cp_elements(655) <= cp_elements(508);
    cp_elements(656) <= cp_elements(525);
    cp_elements(657) <= binary_1514_inst_ack_0;
    binary_1514_inst_req_1 <= cp_elements(657);
    cp_elements(658) <= binary_1514_inst_ack_1;
    array_obj_ref_1518_index_0_resize_req_0 <= cp_elements(658);
    cp_elements(659) <= cp_elements(508);
    cpelement_group_660 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(659) & cp_elements(668));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(660),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1518_final_reg_req_0 <= cp_elements(660);
    cp_elements(661) <= cp_elements(512);
    array_obj_ref_1518_base_resize_req_0 <= cp_elements(661);
    cp_elements(662) <= array_obj_ref_1518_index_0_resize_ack_0;
    array_obj_ref_1518_index_0_rename_req_0 <= cp_elements(662);
    cp_elements(663) <= array_obj_ref_1518_index_0_rename_ack_0;
    array_obj_ref_1518_offset_inst_req_0 <= cp_elements(663);
    cp_elements(664) <= array_obj_ref_1518_offset_inst_ack_0;
    cp_elements(665) <= array_obj_ref_1518_base_resize_ack_0;
    cpelement_group_666 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(664) & cp_elements(665));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(666),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1518_root_address_inst_req_0 <= cp_elements(666);
    cp_elements(667) <= array_obj_ref_1518_root_address_inst_ack_0;
    array_obj_ref_1518_root_address_inst_req_1 <= cp_elements(667);
    cp_elements(668) <= array_obj_ref_1518_root_address_inst_ack_1;
    cp_elements(669) <= array_obj_ref_1518_final_reg_ack_0;
    cpelement_group_670 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(643) & cp_elements(653) & cp_elements(669) & cp_elements(674));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(670),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1521_gather_scatter_req_0 <= cp_elements(670);
    cp_elements(671) <= cp_elements(669);
    ptr_deref_1521_base_resize_req_0 <= cp_elements(671);
    cp_elements(672) <= ptr_deref_1521_base_resize_ack_0;
    ptr_deref_1521_root_address_inst_req_0 <= cp_elements(672);
    cp_elements(673) <= ptr_deref_1521_root_address_inst_ack_0;
    ptr_deref_1521_addr_0_req_0 <= cp_elements(673);
    cp_elements(674) <= ptr_deref_1521_addr_0_ack_0;
    cp_elements(675) <= ptr_deref_1521_gather_scatter_ack_0;
    ptr_deref_1521_store_0_req_0 <= cp_elements(675);
    cp_elements(676) <= ptr_deref_1521_store_0_ack_0;
    cp_elements(677) <= cp_elements(676);
    ptr_deref_1521_store_0_req_1 <= cp_elements(677);
    cp_elements(678) <= ptr_deref_1521_store_0_ack_1;
    cpelement_group_679 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(680) & cp_elements(681));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(679),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1528_inst_req_0 <= cp_elements(679);
    cp_elements(680) <= cp_elements(508);
    cp_elements(681) <= cp_elements(508);
    cp_elements(682) <= binary_1528_inst_ack_0;
    binary_1528_inst_req_1 <= cp_elements(682);
    cp_elements(683) <= binary_1528_inst_ack_1;
    cpelement_group_684 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(683) & cp_elements(685));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(684),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1532_inst_req_0 <= cp_elements(684);
    cp_elements(685) <= cp_elements(508);
    cp_elements(686) <= type_cast_1532_inst_ack_0;
    cpelement_group_687 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(688) & cp_elements(689));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(687),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1538_inst_req_0 <= cp_elements(687);
    cp_elements(688) <= cp_elements(508);
    cp_elements(689) <= cp_elements(525);
    cp_elements(690) <= binary_1538_inst_ack_0;
    binary_1538_inst_req_1 <= cp_elements(690);
    cp_elements(691) <= binary_1538_inst_ack_1;
    array_obj_ref_1542_index_0_resize_req_0 <= cp_elements(691);
    cp_elements(692) <= cp_elements(508);
    cpelement_group_693 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(692) & cp_elements(701));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(693),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1542_final_reg_req_0 <= cp_elements(693);
    cp_elements(694) <= cp_elements(512);
    array_obj_ref_1542_base_resize_req_0 <= cp_elements(694);
    cp_elements(695) <= array_obj_ref_1542_index_0_resize_ack_0;
    array_obj_ref_1542_index_0_rename_req_0 <= cp_elements(695);
    cp_elements(696) <= array_obj_ref_1542_index_0_rename_ack_0;
    array_obj_ref_1542_offset_inst_req_0 <= cp_elements(696);
    cp_elements(697) <= array_obj_ref_1542_offset_inst_ack_0;
    cp_elements(698) <= array_obj_ref_1542_base_resize_ack_0;
    cpelement_group_699 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(697) & cp_elements(698));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(699),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1542_root_address_inst_req_0 <= cp_elements(699);
    cp_elements(700) <= array_obj_ref_1542_root_address_inst_ack_0;
    array_obj_ref_1542_root_address_inst_req_1 <= cp_elements(700);
    cp_elements(701) <= array_obj_ref_1542_root_address_inst_ack_1;
    cp_elements(702) <= array_obj_ref_1542_final_reg_ack_0;
    cpelement_group_703 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(676) & cp_elements(686) & cp_elements(702) & cp_elements(707));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(703),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1545_gather_scatter_req_0 <= cp_elements(703);
    cp_elements(704) <= cp_elements(702);
    ptr_deref_1545_base_resize_req_0 <= cp_elements(704);
    cp_elements(705) <= ptr_deref_1545_base_resize_ack_0;
    ptr_deref_1545_root_address_inst_req_0 <= cp_elements(705);
    cp_elements(706) <= ptr_deref_1545_root_address_inst_ack_0;
    ptr_deref_1545_addr_0_req_0 <= cp_elements(706);
    cp_elements(707) <= ptr_deref_1545_addr_0_ack_0;
    cp_elements(708) <= ptr_deref_1545_gather_scatter_ack_0;
    ptr_deref_1545_store_0_req_0 <= cp_elements(708);
    cp_elements(709) <= ptr_deref_1545_store_0_ack_0;
    cp_elements(710) <= cp_elements(709);
    ptr_deref_1545_store_0_req_1 <= cp_elements(710);
    cp_elements(711) <= ptr_deref_1545_store_0_ack_1;
    cpelement_group_712 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(713) & cp_elements(714));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(712),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1552_inst_req_0 <= cp_elements(712);
    cp_elements(713) <= cp_elements(508);
    cp_elements(714) <= cp_elements(508);
    cp_elements(715) <= binary_1552_inst_ack_0;
    binary_1552_inst_req_1 <= cp_elements(715);
    cp_elements(716) <= binary_1552_inst_ack_1;
    cpelement_group_717 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(716) & cp_elements(718));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(717),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1556_inst_req_0 <= cp_elements(717);
    cp_elements(718) <= cp_elements(508);
    cp_elements(719) <= type_cast_1556_inst_ack_0;
    cpelement_group_720 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(721) & cp_elements(722));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(720),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1562_inst_req_0 <= cp_elements(720);
    cp_elements(721) <= cp_elements(508);
    cp_elements(722) <= cp_elements(525);
    cp_elements(723) <= binary_1562_inst_ack_0;
    binary_1562_inst_req_1 <= cp_elements(723);
    cp_elements(724) <= binary_1562_inst_ack_1;
    array_obj_ref_1566_index_0_resize_req_0 <= cp_elements(724);
    cp_elements(725) <= cp_elements(508);
    cpelement_group_726 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(725) & cp_elements(734));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(726),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1566_final_reg_req_0 <= cp_elements(726);
    cp_elements(727) <= cp_elements(512);
    array_obj_ref_1566_base_resize_req_0 <= cp_elements(727);
    cp_elements(728) <= array_obj_ref_1566_index_0_resize_ack_0;
    array_obj_ref_1566_index_0_rename_req_0 <= cp_elements(728);
    cp_elements(729) <= array_obj_ref_1566_index_0_rename_ack_0;
    array_obj_ref_1566_offset_inst_req_0 <= cp_elements(729);
    cp_elements(730) <= array_obj_ref_1566_offset_inst_ack_0;
    cp_elements(731) <= array_obj_ref_1566_base_resize_ack_0;
    cpelement_group_732 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(730) & cp_elements(731));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(732),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1566_root_address_inst_req_0 <= cp_elements(732);
    cp_elements(733) <= array_obj_ref_1566_root_address_inst_ack_0;
    array_obj_ref_1566_root_address_inst_req_1 <= cp_elements(733);
    cp_elements(734) <= array_obj_ref_1566_root_address_inst_ack_1;
    cp_elements(735) <= array_obj_ref_1566_final_reg_ack_0;
    cpelement_group_736 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(709) & cp_elements(719) & cp_elements(735) & cp_elements(740));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(736),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1569_gather_scatter_req_0 <= cp_elements(736);
    cp_elements(737) <= cp_elements(735);
    ptr_deref_1569_base_resize_req_0 <= cp_elements(737);
    cp_elements(738) <= ptr_deref_1569_base_resize_ack_0;
    ptr_deref_1569_root_address_inst_req_0 <= cp_elements(738);
    cp_elements(739) <= ptr_deref_1569_root_address_inst_ack_0;
    ptr_deref_1569_addr_0_req_0 <= cp_elements(739);
    cp_elements(740) <= ptr_deref_1569_addr_0_ack_0;
    cp_elements(741) <= ptr_deref_1569_gather_scatter_ack_0;
    ptr_deref_1569_store_0_req_0 <= cp_elements(741);
    cp_elements(742) <= ptr_deref_1569_store_0_ack_0;
    cp_elements(743) <= cp_elements(742);
    ptr_deref_1569_store_0_req_1 <= cp_elements(743);
    cp_elements(744) <= ptr_deref_1569_store_0_ack_1;
    cpelement_group_745 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(746) & cp_elements(747));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(745),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1574_inst_req_0 <= cp_elements(745);
    cp_elements(746) <= cp_elements(508);
    cp_elements(747) <= cp_elements(508);
    cp_elements(748) <= type_cast_1574_inst_ack_0;
    cpelement_group_749 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(750) & cp_elements(751));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(749),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1580_inst_req_0 <= cp_elements(749);
    cp_elements(750) <= cp_elements(508);
    cp_elements(751) <= cp_elements(525);
    cp_elements(752) <= binary_1580_inst_ack_0;
    binary_1580_inst_req_1 <= cp_elements(752);
    cp_elements(753) <= binary_1580_inst_ack_1;
    array_obj_ref_1584_index_0_resize_req_0 <= cp_elements(753);
    cp_elements(754) <= cp_elements(508);
    cpelement_group_755 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(754) & cp_elements(763));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(755),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1584_final_reg_req_0 <= cp_elements(755);
    cp_elements(756) <= cp_elements(512);
    array_obj_ref_1584_base_resize_req_0 <= cp_elements(756);
    cp_elements(757) <= array_obj_ref_1584_index_0_resize_ack_0;
    array_obj_ref_1584_index_0_rename_req_0 <= cp_elements(757);
    cp_elements(758) <= array_obj_ref_1584_index_0_rename_ack_0;
    array_obj_ref_1584_offset_inst_req_0 <= cp_elements(758);
    cp_elements(759) <= array_obj_ref_1584_offset_inst_ack_0;
    cp_elements(760) <= array_obj_ref_1584_base_resize_ack_0;
    cpelement_group_761 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(759) & cp_elements(760));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(761),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1584_root_address_inst_req_0 <= cp_elements(761);
    cp_elements(762) <= array_obj_ref_1584_root_address_inst_ack_0;
    array_obj_ref_1584_root_address_inst_req_1 <= cp_elements(762);
    cp_elements(763) <= array_obj_ref_1584_root_address_inst_ack_1;
    cp_elements(764) <= array_obj_ref_1584_final_reg_ack_0;
    cpelement_group_765 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(742) & cp_elements(748) & cp_elements(764) & cp_elements(769));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(765),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1587_gather_scatter_req_0 <= cp_elements(765);
    cp_elements(766) <= cp_elements(764);
    ptr_deref_1587_base_resize_req_0 <= cp_elements(766);
    cp_elements(767) <= ptr_deref_1587_base_resize_ack_0;
    ptr_deref_1587_root_address_inst_req_0 <= cp_elements(767);
    cp_elements(768) <= ptr_deref_1587_root_address_inst_ack_0;
    ptr_deref_1587_addr_0_req_0 <= cp_elements(768);
    cp_elements(769) <= ptr_deref_1587_addr_0_ack_0;
    cp_elements(770) <= ptr_deref_1587_gather_scatter_ack_0;
    ptr_deref_1587_store_0_req_0 <= cp_elements(770);
    cp_elements(771) <= ptr_deref_1587_store_0_ack_0;
    ptr_deref_1587_store_0_req_1 <= cp_elements(771);
    cp_elements(772) <= ptr_deref_1587_store_0_ack_1;
    cpelement_group_773 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(546) & cp_elements(579) & cp_elements(612) & cp_elements(645) & cp_elements(678) & cp_elements(711) & cp_elements(744) & cp_elements(772));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(773),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(774) <= simple_obj_ref_1596_inst_ack_0;
    cp_elements(775) <= OrReduce(cp_elements(2) & cp_elements(35) & cp_elements(774));
    cp_elements(776) <= cp_elements(775);
    simple_obj_ref_981_inst_req_0 <= cp_elements(776);
    cp_elements(777) <= false;
    cp_elements(778) <= cp_elements(777);
    cp_elements(779) <= type_cast_1077_inst_ack_0;
    phi_stmt_1071_req_1 <= cp_elements(779);
    cp_elements(780) <= OrReduce(cp_elements(4) & cp_elements(779));
    cp_elements(781) <= cp_elements(780);
    cp_elements(782) <= phi_stmt_1071_ack_0;
    cp_elements(783) <= OrReduce(cp_elements(5) & cp_elements(7));
    cp_elements(784) <= cp_elements(783);
    simple_obj_ref_1152_inst_req_0 <= cp_elements(784);
    cp_elements(785) <= false;
    cp_elements(786) <= cp_elements(785);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1028_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1028_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1028_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1033_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1033_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1033_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1038_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1038_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1038_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1043_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1043_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1043_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1048_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1057_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1057_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1057_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1062_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1062_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1062_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1067_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1067_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1067_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1093_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1093_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1093_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1093_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1102_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1102_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1102_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1107_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1107_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1107_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1112_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1112_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1112_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1122_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1122_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1122_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1122_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1131_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1131_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1131_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1136_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1136_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1136_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1141_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1141_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1141_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1422_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1422_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1422_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1422_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1446_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1446_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1446_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1446_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1470_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1470_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1470_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1470_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1494_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1494_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1494_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1494_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1518_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1518_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1518_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1518_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1542_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1542_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1542_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1542_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1566_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1566_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1566_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1566_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1584_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1584_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1584_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1584_root_address : std_logic_vector(10 downto 0);
    signal expr_1169_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1169_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_1172_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1172_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal iNsTr_0_967 : std_logic_vector(31 downto 0);
    signal iNsTr_11_1150 : std_logic_vector(31 downto 0);
    signal iNsTr_12_1159 : std_logic_vector(31 downto 0);
    signal iNsTr_22_1595 : std_logic_vector(31 downto 0);
    signal iNsTr_3_980 : std_logic_vector(31 downto 0);
    signal iNsTr_5_990 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1012 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1071 : std_logic_vector(31 downto 0);
    signal ptr_deref_1189_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1189_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1189_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1189_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1189_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1189_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1203_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1203_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1203_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1203_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1203_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1203_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1217_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1217_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1217_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1217_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1217_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1217_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1231_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1231_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1231_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1231_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1231_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1231_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1245_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1245_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1245_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1245_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1245_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1245_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1259_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1259_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1259_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1259_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1259_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1259_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1273_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1273_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1273_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1273_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1273_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1273_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1281_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1281_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1281_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1281_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1281_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1281_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1297_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1297_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1297_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1297_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1297_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1297_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1311_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1311_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1311_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1311_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1311_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1311_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1325_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1325_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1325_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1325_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1325_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1325_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1339_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1339_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1339_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1339_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1339_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1339_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1353_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1353_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1353_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1353_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1353_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1353_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1367_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1367_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1367_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1367_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1367_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1367_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1381_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1381_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1381_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1381_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1381_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1381_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1389_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1389_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1389_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1389_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1389_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1389_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1425_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1425_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1425_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1425_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1425_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1425_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1449_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1449_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1449_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1449_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1449_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1449_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1473_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1473_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1473_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1473_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1473_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1473_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1497_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1497_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1497_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1497_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1497_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1497_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1521_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1521_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1521_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1521_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1521_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1521_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1545_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1545_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1545_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1545_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1545_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1545_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1569_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1569_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1569_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1569_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1569_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1569_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1587_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1587_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1587_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1587_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1587_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1587_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_969_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_969_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_969_word_address_0 : std_logic_vector(3 downto 0);
    signal scevgep147_1123 : std_logic_vector(31 downto 0);
    signal scevgep_1094 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1092_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1092_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1121_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1121_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1421_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1421_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1445_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1445_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1469_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1469_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1493_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1493_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1517_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1517_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1541_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1541_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1565_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1565_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1583_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1583_scaled : std_logic_vector(10 downto 0);
    signal tmp100_1127 : std_logic_vector(31 downto 0);
    signal tmp103_1132 : std_logic_vector(31 downto 0);
    signal tmp106_1137 : std_logic_vector(31 downto 0);
    signal tmp109_1142 : std_logic_vector(31 downto 0);
    signal tmp10_1225 : std_logic_vector(63 downto 0);
    signal tmp110_1397 : std_logic_vector(31 downto 0);
    signal tmp112_1419 : std_logic_vector(31 downto 0);
    signal tmp113_1423 : std_logic_vector(31 downto 0);
    signal tmp115_1443 : std_logic_vector(31 downto 0);
    signal tmp116_1447 : std_logic_vector(31 downto 0);
    signal tmp118_1467 : std_logic_vector(31 downto 0);
    signal tmp119_1471 : std_logic_vector(31 downto 0);
    signal tmp11_1229 : std_logic_vector(7 downto 0);
    signal tmp121_1491 : std_logic_vector(31 downto 0);
    signal tmp122_1495 : std_logic_vector(31 downto 0);
    signal tmp124_1515 : std_logic_vector(31 downto 0);
    signal tmp125_1519 : std_logic_vector(31 downto 0);
    signal tmp127_1539 : std_logic_vector(31 downto 0);
    signal tmp128_1543 : std_logic_vector(31 downto 0);
    signal tmp130_1563 : std_logic_vector(31 downto 0);
    signal tmp131_1567 : std_logic_vector(31 downto 0);
    signal tmp133_1581 : std_logic_vector(31 downto 0);
    signal tmp134_1585 : std_logic_vector(31 downto 0);
    signal tmp138_1090 : std_logic_vector(31 downto 0);
    signal tmp13_1239 : std_logic_vector(63 downto 0);
    signal tmp146_1119 : std_logic_vector(31 downto 0);
    signal tmp14_1243 : std_logic_vector(7 downto 0);
    signal tmp16_1253 : std_logic_vector(63 downto 0);
    signal tmp17_1257 : std_logic_vector(7 downto 0);
    signal tmp19_1267 : std_logic_vector(63 downto 0);
    signal tmp1_1183 : std_logic_vector(63 downto 0);
    signal tmp20_1271 : std_logic_vector(7 downto 0);
    signal tmp22_1279 : std_logic_vector(7 downto 0);
    signal tmp24_1291 : std_logic_vector(63 downto 0);
    signal tmp25_1295 : std_logic_vector(7 downto 0);
    signal tmp27_1305 : std_logic_vector(63 downto 0);
    signal tmp28_1309 : std_logic_vector(7 downto 0);
    signal tmp2_1187 : std_logic_vector(7 downto 0);
    signal tmp2x_xi_999 : std_logic_vector(0 downto 0);
    signal tmp30_1319 : std_logic_vector(63 downto 0);
    signal tmp31_1323 : std_logic_vector(7 downto 0);
    signal tmp33_1333 : std_logic_vector(63 downto 0);
    signal tmp34_1337 : std_logic_vector(7 downto 0);
    signal tmp36_1347 : std_logic_vector(63 downto 0);
    signal tmp37_1351 : std_logic_vector(7 downto 0);
    signal tmp39_1361 : std_logic_vector(63 downto 0);
    signal tmp40_1365 : std_logic_vector(7 downto 0);
    signal tmp42_1375 : std_logic_vector(63 downto 0);
    signal tmp43_1379 : std_logic_vector(7 downto 0);
    signal tmp45_1387 : std_logic_vector(7 downto 0);
    signal tmp47_1409 : std_logic_vector(63 downto 0);
    signal tmp48_1413 : std_logic_vector(7 downto 0);
    signal tmp4_1197 : std_logic_vector(63 downto 0);
    signal tmp4x_xi_1015 : std_logic_vector(31 downto 0);
    signal tmp50_1433 : std_logic_vector(63 downto 0);
    signal tmp51_1437 : std_logic_vector(7 downto 0);
    signal tmp53_1457 : std_logic_vector(63 downto 0);
    signal tmp54_1461 : std_logic_vector(7 downto 0);
    signal tmp56_1481 : std_logic_vector(63 downto 0);
    signal tmp57_1485 : std_logic_vector(7 downto 0);
    signal tmp59_1505 : std_logic_vector(63 downto 0);
    signal tmp5_1201 : std_logic_vector(7 downto 0);
    signal tmp5x_xi_1019 : std_logic_vector(31 downto 0);
    signal tmp60_1509 : std_logic_vector(7 downto 0);
    signal tmp62_1529 : std_logic_vector(63 downto 0);
    signal tmp63_1533 : std_logic_vector(7 downto 0);
    signal tmp65_1553 : std_logic_vector(63 downto 0);
    signal tmp66_1557 : std_logic_vector(7 downto 0);
    signal tmp68_1575 : std_logic_vector(7 downto 0);
    signal tmp70_1024 : std_logic_vector(31 downto 0);
    signal tmp71_1029 : std_logic_vector(31 downto 0);
    signal tmp72_1403 : std_logic_vector(31 downto 0);
    signal tmp74_1153 : std_logic_vector(63 downto 0);
    signal tmp75_1162 : std_logic_vector(7 downto 0);
    signal tmp76_1166 : std_logic_vector(31 downto 0);
    signal tmp78_1034 : std_logic_vector(31 downto 0);
    signal tmp79_1039 : std_logic_vector(31 downto 0);
    signal tmp7_1211 : std_logic_vector(63 downto 0);
    signal tmp80_1044 : std_logic_vector(31 downto 0);
    signal tmp81_1049 : std_logic_vector(31 downto 0);
    signal tmp82_1053 : std_logic_vector(31 downto 0);
    signal tmp83_1058 : std_logic_vector(31 downto 0);
    signal tmp84_1063 : std_logic_vector(31 downto 0);
    signal tmp85_1068 : std_logic_vector(31 downto 0);
    signal tmp88_1098 : std_logic_vector(31 downto 0);
    signal tmp8_1215 : std_logic_vector(7 downto 0);
    signal tmp91_1103 : std_logic_vector(31 downto 0);
    signal tmp94_1108 : std_logic_vector(31 downto 0);
    signal tmp97_1113 : std_logic_vector(31 downto 0);
    signal tmp_1084 : std_logic_vector(31 downto 0);
    signal tmpx_xi_993 : std_logic_vector(7 downto 0);
    signal type_cast_1075_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1077_wire : std_logic_vector(31 downto 0);
    signal type_cast_1082_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1088_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1117_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1181_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1195_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1209_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1223_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1237_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1251_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1265_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1289_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1303_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1317_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1331_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1345_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1359_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1373_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1395_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1407_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1417_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1431_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1441_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1455_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1465_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1479_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1489_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1503_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1527_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1537_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1551_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1561_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1579_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_971_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_983_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1028_final_offset <= "00000001000";
    array_obj_ref_1033_final_offset <= "00000000001";
    array_obj_ref_1038_final_offset <= "00000000010";
    array_obj_ref_1043_final_offset <= "00000000011";
    array_obj_ref_1048_final_offset <= "00000000100";
    array_obj_ref_1057_final_offset <= "00000000101";
    array_obj_ref_1062_final_offset <= "00000000110";
    array_obj_ref_1067_final_offset <= "00000000111";
    array_obj_ref_1093_offset_scale_factor_0 <= "00000000100";
    array_obj_ref_1102_final_offset <= "00000000001";
    array_obj_ref_1107_final_offset <= "00000000010";
    array_obj_ref_1112_final_offset <= "00000000011";
    array_obj_ref_1122_offset_scale_factor_0 <= "00000000100";
    array_obj_ref_1131_final_offset <= "00000000001";
    array_obj_ref_1136_final_offset <= "00000000010";
    array_obj_ref_1141_final_offset <= "00000000011";
    array_obj_ref_1422_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1446_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1470_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1494_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1518_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1542_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1566_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1584_offset_scale_factor_0 <= "00000000001";
    expr_1169_wire_constant <= "00000000000000000000000011111111";
    expr_1172_wire_constant <= "00000000000000000000000000000000";
    iNsTr_0_967 <= "00000000000000000000000000000000";
    iNsTr_11_1150 <= "00000000000000000000000000000000";
    iNsTr_12_1159 <= "00000000000000000000000000000000";
    iNsTr_22_1595 <= "00000000000000000000000000000000";
    iNsTr_3_980 <= "00000000000000000000000000000000";
    iNsTr_5_990 <= "00000000000000000000000000000000";
    iNsTr_7_1012 <= "00000000000000000000000000000000";
    ptr_deref_1189_word_offset_0 <= "00000000000";
    ptr_deref_1203_word_offset_0 <= "00000000000";
    ptr_deref_1217_word_offset_0 <= "00000000000";
    ptr_deref_1231_word_offset_0 <= "00000000000";
    ptr_deref_1245_word_offset_0 <= "00000000000";
    ptr_deref_1259_word_offset_0 <= "00000000000";
    ptr_deref_1273_word_offset_0 <= "00000000000";
    ptr_deref_1281_word_offset_0 <= "00000000000";
    ptr_deref_1297_word_offset_0 <= "00000000000";
    ptr_deref_1311_word_offset_0 <= "00000000000";
    ptr_deref_1325_word_offset_0 <= "00000000000";
    ptr_deref_1339_word_offset_0 <= "00000000000";
    ptr_deref_1353_word_offset_0 <= "00000000000";
    ptr_deref_1367_word_offset_0 <= "00000000000";
    ptr_deref_1381_word_offset_0 <= "00000000000";
    ptr_deref_1389_word_offset_0 <= "00000000000";
    ptr_deref_1425_word_offset_0 <= "00000000000";
    ptr_deref_1449_word_offset_0 <= "00000000000";
    ptr_deref_1473_word_offset_0 <= "00000000000";
    ptr_deref_1497_word_offset_0 <= "00000000000";
    ptr_deref_1521_word_offset_0 <= "00000000000";
    ptr_deref_1545_word_offset_0 <= "00000000000";
    ptr_deref_1569_word_offset_0 <= "00000000000";
    ptr_deref_1587_word_offset_0 <= "00000000000";
    ptr_deref_969_word_address_0 <= "0000";
    type_cast_1075_wire_constant <= "00000000000000000000000000000000";
    type_cast_1082_wire_constant <= "00000000000000000000000000000001";
    type_cast_1088_wire_constant <= "00000000000000000000000000000010";
    type_cast_1117_wire_constant <= "00000000000000000000000000000011";
    type_cast_1181_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1209_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1223_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1237_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1251_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1265_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1289_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1303_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1317_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1331_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1345_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1359_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1373_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1395_wire_constant <= "00000000000000000000000000000001";
    type_cast_1407_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1417_wire_constant <= "00000000000000000000000000000011";
    type_cast_1431_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1441_wire_constant <= "00000000000000000000000000000001";
    type_cast_1455_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1465_wire_constant <= "00000000000000000000000000000010";
    type_cast_1479_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1489_wire_constant <= "00000000000000000000000000000011";
    type_cast_1503_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1513_wire_constant <= "00000000000000000000000000000100";
    type_cast_1527_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1537_wire_constant <= "00000000000000000000000000000101";
    type_cast_1551_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1561_wire_constant <= "00000000000000000000000000000110";
    type_cast_1579_wire_constant <= "00000000000000000000000000000111";
    type_cast_971_wire_constant <= "00000001";
    type_cast_983_wire_constant <= "00000010";
    type_cast_997_wire_constant <= "00000011";
    phi_stmt_1071: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1075_wire_constant & type_cast_1077_wire;
      req <= phi_stmt_1071_req_0 & phi_stmt_1071_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1071_ack_0,
          idata => idata,
          odata => iNsTr_9_1071,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1071
    array_obj_ref_1028_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp5x_xi_1019, dout => array_obj_ref_1028_resized_base_address, req => array_obj_ref_1028_base_resize_req_0, ack => array_obj_ref_1028_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1028_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1028_root_address, dout => tmp71_1029, req => array_obj_ref_1028_final_reg_req_0, ack => array_obj_ref_1028_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1033_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1024, dout => array_obj_ref_1033_resized_base_address, req => array_obj_ref_1033_base_resize_req_0, ack => array_obj_ref_1033_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1033_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1033_root_address, dout => tmp78_1034, req => array_obj_ref_1033_final_reg_req_0, ack => array_obj_ref_1033_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1038_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1024, dout => array_obj_ref_1038_resized_base_address, req => array_obj_ref_1038_base_resize_req_0, ack => array_obj_ref_1038_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1038_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1038_root_address, dout => tmp79_1039, req => array_obj_ref_1038_final_reg_req_0, ack => array_obj_ref_1038_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1043_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1024, dout => array_obj_ref_1043_resized_base_address, req => array_obj_ref_1043_base_resize_req_0, ack => array_obj_ref_1043_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1043_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1043_root_address, dout => tmp80_1044, req => array_obj_ref_1043_final_reg_req_0, ack => array_obj_ref_1043_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1048_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp5x_xi_1019, dout => array_obj_ref_1048_resized_base_address, req => array_obj_ref_1048_base_resize_req_0, ack => array_obj_ref_1048_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1048_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1048_root_address, dout => tmp81_1049, req => array_obj_ref_1048_final_reg_req_0, ack => array_obj_ref_1048_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1057_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1024, dout => array_obj_ref_1057_resized_base_address, req => array_obj_ref_1057_base_resize_req_0, ack => array_obj_ref_1057_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1057_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1057_root_address, dout => tmp83_1058, req => array_obj_ref_1057_final_reg_req_0, ack => array_obj_ref_1057_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1062_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1024, dout => array_obj_ref_1062_resized_base_address, req => array_obj_ref_1062_base_resize_req_0, ack => array_obj_ref_1062_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1062_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1062_root_address, dout => tmp84_1063, req => array_obj_ref_1062_final_reg_req_0, ack => array_obj_ref_1062_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1067_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1024, dout => array_obj_ref_1067_resized_base_address, req => array_obj_ref_1067_base_resize_req_0, ack => array_obj_ref_1067_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1067_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1067_root_address, dout => tmp85_1068, req => array_obj_ref_1067_final_reg_req_0, ack => array_obj_ref_1067_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1093_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp5x_xi_1019, dout => array_obj_ref_1093_resized_base_address, req => array_obj_ref_1093_base_resize_req_0, ack => array_obj_ref_1093_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1093_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1093_root_address, dout => scevgep_1094, req => array_obj_ref_1093_final_reg_req_0, ack => array_obj_ref_1093_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1093_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp138_1090, dout => simple_obj_ref_1092_resized, req => array_obj_ref_1093_index_0_resize_req_0, ack => array_obj_ref_1093_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1093_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1092_scaled, dout => array_obj_ref_1093_final_offset, req => array_obj_ref_1093_offset_inst_req_0, ack => array_obj_ref_1093_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1102_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp88_1098, dout => array_obj_ref_1102_resized_base_address, req => array_obj_ref_1102_base_resize_req_0, ack => array_obj_ref_1102_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1102_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1102_root_address, dout => tmp91_1103, req => array_obj_ref_1102_final_reg_req_0, ack => array_obj_ref_1102_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1107_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp88_1098, dout => array_obj_ref_1107_resized_base_address, req => array_obj_ref_1107_base_resize_req_0, ack => array_obj_ref_1107_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1107_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1107_root_address, dout => tmp94_1108, req => array_obj_ref_1107_final_reg_req_0, ack => array_obj_ref_1107_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1112_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp88_1098, dout => array_obj_ref_1112_resized_base_address, req => array_obj_ref_1112_base_resize_req_0, ack => array_obj_ref_1112_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1112_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1112_root_address, dout => tmp97_1113, req => array_obj_ref_1112_final_reg_req_0, ack => array_obj_ref_1112_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1122_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp5x_xi_1019, dout => array_obj_ref_1122_resized_base_address, req => array_obj_ref_1122_base_resize_req_0, ack => array_obj_ref_1122_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1122_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1122_root_address, dout => scevgep147_1123, req => array_obj_ref_1122_final_reg_req_0, ack => array_obj_ref_1122_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1122_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp146_1119, dout => simple_obj_ref_1121_resized, req => array_obj_ref_1122_index_0_resize_req_0, ack => array_obj_ref_1122_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1122_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1121_scaled, dout => array_obj_ref_1122_final_offset, req => array_obj_ref_1122_offset_inst_req_0, ack => array_obj_ref_1122_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1131_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp100_1127, dout => array_obj_ref_1131_resized_base_address, req => array_obj_ref_1131_base_resize_req_0, ack => array_obj_ref_1131_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1131_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1131_root_address, dout => tmp103_1132, req => array_obj_ref_1131_final_reg_req_0, ack => array_obj_ref_1131_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1136_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp100_1127, dout => array_obj_ref_1136_resized_base_address, req => array_obj_ref_1136_base_resize_req_0, ack => array_obj_ref_1136_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1136_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1136_root_address, dout => tmp106_1137, req => array_obj_ref_1136_final_reg_req_0, ack => array_obj_ref_1136_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1141_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp100_1127, dout => array_obj_ref_1141_resized_base_address, req => array_obj_ref_1141_base_resize_req_0, ack => array_obj_ref_1141_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1141_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1141_root_address, dout => tmp109_1142, req => array_obj_ref_1141_final_reg_req_0, ack => array_obj_ref_1141_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1422_resized_base_address, req => array_obj_ref_1422_base_resize_req_0, ack => array_obj_ref_1422_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1422_root_address, dout => tmp113_1423, req => array_obj_ref_1422_final_reg_req_0, ack => array_obj_ref_1422_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp112_1419, dout => simple_obj_ref_1421_resized, req => array_obj_ref_1422_index_0_resize_req_0, ack => array_obj_ref_1422_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1421_scaled, dout => array_obj_ref_1422_final_offset, req => array_obj_ref_1422_offset_inst_req_0, ack => array_obj_ref_1422_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1446_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1446_resized_base_address, req => array_obj_ref_1446_base_resize_req_0, ack => array_obj_ref_1446_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1446_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1446_root_address, dout => tmp116_1447, req => array_obj_ref_1446_final_reg_req_0, ack => array_obj_ref_1446_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1446_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp115_1443, dout => simple_obj_ref_1445_resized, req => array_obj_ref_1446_index_0_resize_req_0, ack => array_obj_ref_1446_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1446_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1445_scaled, dout => array_obj_ref_1446_final_offset, req => array_obj_ref_1446_offset_inst_req_0, ack => array_obj_ref_1446_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1470_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1470_resized_base_address, req => array_obj_ref_1470_base_resize_req_0, ack => array_obj_ref_1470_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1470_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1470_root_address, dout => tmp119_1471, req => array_obj_ref_1470_final_reg_req_0, ack => array_obj_ref_1470_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1470_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp118_1467, dout => simple_obj_ref_1469_resized, req => array_obj_ref_1470_index_0_resize_req_0, ack => array_obj_ref_1470_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1470_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1469_scaled, dout => array_obj_ref_1470_final_offset, req => array_obj_ref_1470_offset_inst_req_0, ack => array_obj_ref_1470_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1494_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1494_resized_base_address, req => array_obj_ref_1494_base_resize_req_0, ack => array_obj_ref_1494_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1494_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1494_root_address, dout => tmp122_1495, req => array_obj_ref_1494_final_reg_req_0, ack => array_obj_ref_1494_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1494_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp121_1491, dout => simple_obj_ref_1493_resized, req => array_obj_ref_1494_index_0_resize_req_0, ack => array_obj_ref_1494_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1494_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1493_scaled, dout => array_obj_ref_1494_final_offset, req => array_obj_ref_1494_offset_inst_req_0, ack => array_obj_ref_1494_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1518_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1518_resized_base_address, req => array_obj_ref_1518_base_resize_req_0, ack => array_obj_ref_1518_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1518_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1518_root_address, dout => tmp125_1519, req => array_obj_ref_1518_final_reg_req_0, ack => array_obj_ref_1518_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1518_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1515, dout => simple_obj_ref_1517_resized, req => array_obj_ref_1518_index_0_resize_req_0, ack => array_obj_ref_1518_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1518_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1517_scaled, dout => array_obj_ref_1518_final_offset, req => array_obj_ref_1518_offset_inst_req_0, ack => array_obj_ref_1518_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1542_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1542_resized_base_address, req => array_obj_ref_1542_base_resize_req_0, ack => array_obj_ref_1542_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1542_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1542_root_address, dout => tmp128_1543, req => array_obj_ref_1542_final_reg_req_0, ack => array_obj_ref_1542_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1542_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp127_1539, dout => simple_obj_ref_1541_resized, req => array_obj_ref_1542_index_0_resize_req_0, ack => array_obj_ref_1542_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1542_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1541_scaled, dout => array_obj_ref_1542_final_offset, req => array_obj_ref_1542_offset_inst_req_0, ack => array_obj_ref_1542_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1566_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1566_resized_base_address, req => array_obj_ref_1566_base_resize_req_0, ack => array_obj_ref_1566_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1566_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1566_root_address, dout => tmp131_1567, req => array_obj_ref_1566_final_reg_req_0, ack => array_obj_ref_1566_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1566_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp130_1563, dout => simple_obj_ref_1565_resized, req => array_obj_ref_1566_index_0_resize_req_0, ack => array_obj_ref_1566_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1566_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1565_scaled, dout => array_obj_ref_1566_final_offset, req => array_obj_ref_1566_offset_inst_req_0, ack => array_obj_ref_1566_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1584_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp72_1403, dout => array_obj_ref_1584_resized_base_address, req => array_obj_ref_1584_base_resize_req_0, ack => array_obj_ref_1584_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1584_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1584_root_address, dout => tmp134_1585, req => array_obj_ref_1584_final_reg_req_0, ack => array_obj_ref_1584_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1584_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp133_1581, dout => simple_obj_ref_1583_resized, req => array_obj_ref_1584_index_0_resize_req_0, ack => array_obj_ref_1584_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1584_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1583_scaled, dout => array_obj_ref_1584_final_offset, req => array_obj_ref_1584_offset_inst_req_0, ack => array_obj_ref_1584_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1189_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1024, dout => ptr_deref_1189_resized_base_address, req => ptr_deref_1189_base_resize_req_0, ack => ptr_deref_1189_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1203_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp78_1034, dout => ptr_deref_1203_resized_base_address, req => ptr_deref_1203_base_resize_req_0, ack => ptr_deref_1203_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1217_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp79_1039, dout => ptr_deref_1217_resized_base_address, req => ptr_deref_1217_base_resize_req_0, ack => ptr_deref_1217_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1231_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp80_1044, dout => ptr_deref_1231_resized_base_address, req => ptr_deref_1231_base_resize_req_0, ack => ptr_deref_1231_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1245_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp82_1053, dout => ptr_deref_1245_resized_base_address, req => ptr_deref_1245_base_resize_req_0, ack => ptr_deref_1245_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1259_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp83_1058, dout => ptr_deref_1259_resized_base_address, req => ptr_deref_1259_base_resize_req_0, ack => ptr_deref_1259_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1273_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp84_1063, dout => ptr_deref_1273_resized_base_address, req => ptr_deref_1273_base_resize_req_0, ack => ptr_deref_1273_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1281_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp85_1068, dout => ptr_deref_1281_resized_base_address, req => ptr_deref_1281_base_resize_req_0, ack => ptr_deref_1281_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1297_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp88_1098, dout => ptr_deref_1297_resized_base_address, req => ptr_deref_1297_base_resize_req_0, ack => ptr_deref_1297_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1311_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp91_1103, dout => ptr_deref_1311_resized_base_address, req => ptr_deref_1311_base_resize_req_0, ack => ptr_deref_1311_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1325_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp94_1108, dout => ptr_deref_1325_resized_base_address, req => ptr_deref_1325_base_resize_req_0, ack => ptr_deref_1325_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1339_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp97_1113, dout => ptr_deref_1339_resized_base_address, req => ptr_deref_1339_base_resize_req_0, ack => ptr_deref_1339_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1353_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp100_1127, dout => ptr_deref_1353_resized_base_address, req => ptr_deref_1353_base_resize_req_0, ack => ptr_deref_1353_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1367_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp103_1132, dout => ptr_deref_1367_resized_base_address, req => ptr_deref_1367_base_resize_req_0, ack => ptr_deref_1367_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1381_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp106_1137, dout => ptr_deref_1381_resized_base_address, req => ptr_deref_1381_base_resize_req_0, ack => ptr_deref_1381_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1389_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp109_1142, dout => ptr_deref_1389_resized_base_address, req => ptr_deref_1389_base_resize_req_0, ack => ptr_deref_1389_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1425_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp113_1423, dout => ptr_deref_1425_resized_base_address, req => ptr_deref_1425_base_resize_req_0, ack => ptr_deref_1425_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1449_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp116_1447, dout => ptr_deref_1449_resized_base_address, req => ptr_deref_1449_base_resize_req_0, ack => ptr_deref_1449_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1473_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp119_1471, dout => ptr_deref_1473_resized_base_address, req => ptr_deref_1473_base_resize_req_0, ack => ptr_deref_1473_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1497_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp122_1495, dout => ptr_deref_1497_resized_base_address, req => ptr_deref_1497_base_resize_req_0, ack => ptr_deref_1497_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1521_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_1519, dout => ptr_deref_1521_resized_base_address, req => ptr_deref_1521_base_resize_req_0, ack => ptr_deref_1521_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1545_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp128_1543, dout => ptr_deref_1545_resized_base_address, req => ptr_deref_1545_base_resize_req_0, ack => ptr_deref_1545_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1569_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp131_1567, dout => ptr_deref_1569_resized_base_address, req => ptr_deref_1569_base_resize_req_0, ack => ptr_deref_1569_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1587_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp134_1585, dout => ptr_deref_1587_resized_base_address, req => ptr_deref_1587_base_resize_req_0, ack => ptr_deref_1587_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1018_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp4x_xi_1015, dout => tmp5x_xi_1019, req => type_cast_1018_inst_req_0, ack => type_cast_1018_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1023_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp4x_xi_1015, dout => tmp70_1024, req => type_cast_1023_inst_req_0, ack => type_cast_1023_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1052_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp81_1049, dout => tmp82_1053, req => type_cast_1052_inst_req_0, ack => type_cast_1052_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1077_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp110_1397, dout => type_cast_1077_wire, req => type_cast_1077_inst_req_0, ack => type_cast_1077_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1097_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => scevgep_1094, dout => tmp88_1098, req => type_cast_1097_inst_req_0, ack => type_cast_1097_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1126_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => scevgep147_1123, dout => tmp100_1127, req => type_cast_1126_inst_req_0, ack => type_cast_1126_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1165_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 32, flow_through => false ) 
      port map( din => tmp75_1162, dout => tmp76_1166, req => type_cast_1165_inst_req_0, ack => type_cast_1165_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1186_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp1_1183, dout => tmp2_1187, req => type_cast_1186_inst_req_0, ack => type_cast_1186_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1200_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp4_1197, dout => tmp5_1201, req => type_cast_1200_inst_req_0, ack => type_cast_1200_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1214_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp7_1211, dout => tmp8_1215, req => type_cast_1214_inst_req_0, ack => type_cast_1214_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1228_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp10_1225, dout => tmp11_1229, req => type_cast_1228_inst_req_0, ack => type_cast_1228_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1242_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp13_1239, dout => tmp14_1243, req => type_cast_1242_inst_req_0, ack => type_cast_1242_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1256_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp16_1253, dout => tmp17_1257, req => type_cast_1256_inst_req_0, ack => type_cast_1256_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1270_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp19_1267, dout => tmp20_1271, req => type_cast_1270_inst_req_0, ack => type_cast_1270_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1278_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp74_1153, dout => tmp22_1279, req => type_cast_1278_inst_req_0, ack => type_cast_1278_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1294_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp24_1291, dout => tmp25_1295, req => type_cast_1294_inst_req_0, ack => type_cast_1294_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1308_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp27_1305, dout => tmp28_1309, req => type_cast_1308_inst_req_0, ack => type_cast_1308_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1322_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp30_1319, dout => tmp31_1323, req => type_cast_1322_inst_req_0, ack => type_cast_1322_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1336_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp33_1333, dout => tmp34_1337, req => type_cast_1336_inst_req_0, ack => type_cast_1336_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1350_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp36_1347, dout => tmp37_1351, req => type_cast_1350_inst_req_0, ack => type_cast_1350_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1364_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp39_1361, dout => tmp40_1365, req => type_cast_1364_inst_req_0, ack => type_cast_1364_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1378_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp42_1375, dout => tmp43_1379, req => type_cast_1378_inst_req_0, ack => type_cast_1378_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1386_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp74_1153, dout => tmp45_1387, req => type_cast_1386_inst_req_0, ack => type_cast_1386_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1402_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp71_1029, dout => tmp72_1403, req => type_cast_1402_inst_req_0, ack => type_cast_1402_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1412_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp47_1409, dout => tmp48_1413, req => type_cast_1412_inst_req_0, ack => type_cast_1412_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1436_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp50_1433, dout => tmp51_1437, req => type_cast_1436_inst_req_0, ack => type_cast_1436_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1460_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp53_1457, dout => tmp54_1461, req => type_cast_1460_inst_req_0, ack => type_cast_1460_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1484_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp56_1481, dout => tmp57_1485, req => type_cast_1484_inst_req_0, ack => type_cast_1484_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1508_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp59_1505, dout => tmp60_1509, req => type_cast_1508_inst_req_0, ack => type_cast_1508_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1532_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp62_1529, dout => tmp63_1533, req => type_cast_1532_inst_req_0, ack => type_cast_1532_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1556_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp65_1553, dout => tmp66_1557, req => type_cast_1556_inst_req_0, ack => type_cast_1556_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1574_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp74_1153, dout => tmp68_1575, req => type_cast_1574_inst_req_0, ack => type_cast_1574_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1422_index_0_rename_ack_0 <= array_obj_ref_1422_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1421_resized;
      simple_obj_ref_1421_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1446_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1446_index_0_rename_ack_0 <= array_obj_ref_1446_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1445_resized;
      simple_obj_ref_1445_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1470_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1470_index_0_rename_ack_0 <= array_obj_ref_1470_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1469_resized;
      simple_obj_ref_1469_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1494_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1494_index_0_rename_ack_0 <= array_obj_ref_1494_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1493_resized;
      simple_obj_ref_1493_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1518_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1518_index_0_rename_ack_0 <= array_obj_ref_1518_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1517_resized;
      simple_obj_ref_1517_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1542_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1542_index_0_rename_ack_0 <= array_obj_ref_1542_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1541_resized;
      simple_obj_ref_1541_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1566_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1566_index_0_rename_ack_0 <= array_obj_ref_1566_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1565_resized;
      simple_obj_ref_1565_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1584_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1584_index_0_rename_ack_0 <= array_obj_ref_1584_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1583_resized;
      simple_obj_ref_1583_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1189_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1189_addr_0_ack_0 <= ptr_deref_1189_addr_0_req_0;
      aggregated_sig <= ptr_deref_1189_root_address;
      ptr_deref_1189_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1189_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1189_gather_scatter_ack_0 <= ptr_deref_1189_gather_scatter_req_0;
      aggregated_sig <= tmp2_1187;
      ptr_deref_1189_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1189_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1189_root_address_inst_ack_0 <= ptr_deref_1189_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1189_resized_base_address;
      ptr_deref_1189_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1203_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1203_addr_0_ack_0 <= ptr_deref_1203_addr_0_req_0;
      aggregated_sig <= ptr_deref_1203_root_address;
      ptr_deref_1203_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1203_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1203_gather_scatter_ack_0 <= ptr_deref_1203_gather_scatter_req_0;
      aggregated_sig <= tmp5_1201;
      ptr_deref_1203_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1203_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1203_root_address_inst_ack_0 <= ptr_deref_1203_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1203_resized_base_address;
      ptr_deref_1203_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1217_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1217_addr_0_ack_0 <= ptr_deref_1217_addr_0_req_0;
      aggregated_sig <= ptr_deref_1217_root_address;
      ptr_deref_1217_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1217_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1217_gather_scatter_ack_0 <= ptr_deref_1217_gather_scatter_req_0;
      aggregated_sig <= tmp8_1215;
      ptr_deref_1217_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1217_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1217_root_address_inst_ack_0 <= ptr_deref_1217_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1217_resized_base_address;
      ptr_deref_1217_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1231_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1231_addr_0_ack_0 <= ptr_deref_1231_addr_0_req_0;
      aggregated_sig <= ptr_deref_1231_root_address;
      ptr_deref_1231_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1231_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1231_gather_scatter_ack_0 <= ptr_deref_1231_gather_scatter_req_0;
      aggregated_sig <= tmp11_1229;
      ptr_deref_1231_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1231_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1231_root_address_inst_ack_0 <= ptr_deref_1231_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1231_resized_base_address;
      ptr_deref_1231_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1245_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1245_addr_0_ack_0 <= ptr_deref_1245_addr_0_req_0;
      aggregated_sig <= ptr_deref_1245_root_address;
      ptr_deref_1245_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1245_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1245_gather_scatter_ack_0 <= ptr_deref_1245_gather_scatter_req_0;
      aggregated_sig <= tmp14_1243;
      ptr_deref_1245_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1245_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1245_root_address_inst_ack_0 <= ptr_deref_1245_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1245_resized_base_address;
      ptr_deref_1245_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1259_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1259_addr_0_ack_0 <= ptr_deref_1259_addr_0_req_0;
      aggregated_sig <= ptr_deref_1259_root_address;
      ptr_deref_1259_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1259_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1259_gather_scatter_ack_0 <= ptr_deref_1259_gather_scatter_req_0;
      aggregated_sig <= tmp17_1257;
      ptr_deref_1259_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1259_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1259_root_address_inst_ack_0 <= ptr_deref_1259_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1259_resized_base_address;
      ptr_deref_1259_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1273_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1273_addr_0_ack_0 <= ptr_deref_1273_addr_0_req_0;
      aggregated_sig <= ptr_deref_1273_root_address;
      ptr_deref_1273_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1273_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1273_gather_scatter_ack_0 <= ptr_deref_1273_gather_scatter_req_0;
      aggregated_sig <= tmp20_1271;
      ptr_deref_1273_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1273_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1273_root_address_inst_ack_0 <= ptr_deref_1273_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1273_resized_base_address;
      ptr_deref_1273_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1281_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1281_addr_0_ack_0 <= ptr_deref_1281_addr_0_req_0;
      aggregated_sig <= ptr_deref_1281_root_address;
      ptr_deref_1281_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1281_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1281_gather_scatter_ack_0 <= ptr_deref_1281_gather_scatter_req_0;
      aggregated_sig <= tmp22_1279;
      ptr_deref_1281_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1281_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1281_root_address_inst_ack_0 <= ptr_deref_1281_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1281_resized_base_address;
      ptr_deref_1281_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1297_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1297_addr_0_ack_0 <= ptr_deref_1297_addr_0_req_0;
      aggregated_sig <= ptr_deref_1297_root_address;
      ptr_deref_1297_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1297_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1297_gather_scatter_ack_0 <= ptr_deref_1297_gather_scatter_req_0;
      aggregated_sig <= tmp25_1295;
      ptr_deref_1297_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1297_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1297_root_address_inst_ack_0 <= ptr_deref_1297_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1297_resized_base_address;
      ptr_deref_1297_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1311_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1311_addr_0_ack_0 <= ptr_deref_1311_addr_0_req_0;
      aggregated_sig <= ptr_deref_1311_root_address;
      ptr_deref_1311_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1311_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1311_gather_scatter_ack_0 <= ptr_deref_1311_gather_scatter_req_0;
      aggregated_sig <= tmp28_1309;
      ptr_deref_1311_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1311_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1311_root_address_inst_ack_0 <= ptr_deref_1311_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1311_resized_base_address;
      ptr_deref_1311_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1325_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1325_addr_0_ack_0 <= ptr_deref_1325_addr_0_req_0;
      aggregated_sig <= ptr_deref_1325_root_address;
      ptr_deref_1325_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1325_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1325_gather_scatter_ack_0 <= ptr_deref_1325_gather_scatter_req_0;
      aggregated_sig <= tmp31_1323;
      ptr_deref_1325_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1325_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1325_root_address_inst_ack_0 <= ptr_deref_1325_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1325_resized_base_address;
      ptr_deref_1325_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1339_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1339_addr_0_ack_0 <= ptr_deref_1339_addr_0_req_0;
      aggregated_sig <= ptr_deref_1339_root_address;
      ptr_deref_1339_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1339_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1339_gather_scatter_ack_0 <= ptr_deref_1339_gather_scatter_req_0;
      aggregated_sig <= tmp34_1337;
      ptr_deref_1339_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1339_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1339_root_address_inst_ack_0 <= ptr_deref_1339_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1339_resized_base_address;
      ptr_deref_1339_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1353_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1353_addr_0_ack_0 <= ptr_deref_1353_addr_0_req_0;
      aggregated_sig <= ptr_deref_1353_root_address;
      ptr_deref_1353_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1353_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1353_gather_scatter_ack_0 <= ptr_deref_1353_gather_scatter_req_0;
      aggregated_sig <= tmp37_1351;
      ptr_deref_1353_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1353_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1353_root_address_inst_ack_0 <= ptr_deref_1353_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1353_resized_base_address;
      ptr_deref_1353_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1367_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1367_addr_0_ack_0 <= ptr_deref_1367_addr_0_req_0;
      aggregated_sig <= ptr_deref_1367_root_address;
      ptr_deref_1367_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1367_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1367_gather_scatter_ack_0 <= ptr_deref_1367_gather_scatter_req_0;
      aggregated_sig <= tmp40_1365;
      ptr_deref_1367_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1367_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1367_root_address_inst_ack_0 <= ptr_deref_1367_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1367_resized_base_address;
      ptr_deref_1367_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1381_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1381_addr_0_ack_0 <= ptr_deref_1381_addr_0_req_0;
      aggregated_sig <= ptr_deref_1381_root_address;
      ptr_deref_1381_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1381_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1381_gather_scatter_ack_0 <= ptr_deref_1381_gather_scatter_req_0;
      aggregated_sig <= tmp43_1379;
      ptr_deref_1381_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1381_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1381_root_address_inst_ack_0 <= ptr_deref_1381_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1381_resized_base_address;
      ptr_deref_1381_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1389_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1389_addr_0_ack_0 <= ptr_deref_1389_addr_0_req_0;
      aggregated_sig <= ptr_deref_1389_root_address;
      ptr_deref_1389_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1389_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1389_gather_scatter_ack_0 <= ptr_deref_1389_gather_scatter_req_0;
      aggregated_sig <= tmp45_1387;
      ptr_deref_1389_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1389_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1389_root_address_inst_ack_0 <= ptr_deref_1389_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1389_resized_base_address;
      ptr_deref_1389_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1425_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1425_addr_0_ack_0 <= ptr_deref_1425_addr_0_req_0;
      aggregated_sig <= ptr_deref_1425_root_address;
      ptr_deref_1425_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1425_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1425_gather_scatter_ack_0 <= ptr_deref_1425_gather_scatter_req_0;
      aggregated_sig <= tmp48_1413;
      ptr_deref_1425_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1425_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1425_root_address_inst_ack_0 <= ptr_deref_1425_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1425_resized_base_address;
      ptr_deref_1425_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1449_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1449_addr_0_ack_0 <= ptr_deref_1449_addr_0_req_0;
      aggregated_sig <= ptr_deref_1449_root_address;
      ptr_deref_1449_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1449_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1449_gather_scatter_ack_0 <= ptr_deref_1449_gather_scatter_req_0;
      aggregated_sig <= tmp51_1437;
      ptr_deref_1449_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1449_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1449_root_address_inst_ack_0 <= ptr_deref_1449_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1449_resized_base_address;
      ptr_deref_1449_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1473_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1473_addr_0_ack_0 <= ptr_deref_1473_addr_0_req_0;
      aggregated_sig <= ptr_deref_1473_root_address;
      ptr_deref_1473_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1473_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1473_gather_scatter_ack_0 <= ptr_deref_1473_gather_scatter_req_0;
      aggregated_sig <= tmp54_1461;
      ptr_deref_1473_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1473_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1473_root_address_inst_ack_0 <= ptr_deref_1473_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1473_resized_base_address;
      ptr_deref_1473_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1497_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1497_addr_0_ack_0 <= ptr_deref_1497_addr_0_req_0;
      aggregated_sig <= ptr_deref_1497_root_address;
      ptr_deref_1497_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1497_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1497_gather_scatter_ack_0 <= ptr_deref_1497_gather_scatter_req_0;
      aggregated_sig <= tmp57_1485;
      ptr_deref_1497_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1497_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1497_root_address_inst_ack_0 <= ptr_deref_1497_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1497_resized_base_address;
      ptr_deref_1497_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1521_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1521_addr_0_ack_0 <= ptr_deref_1521_addr_0_req_0;
      aggregated_sig <= ptr_deref_1521_root_address;
      ptr_deref_1521_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1521_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1521_gather_scatter_ack_0 <= ptr_deref_1521_gather_scatter_req_0;
      aggregated_sig <= tmp60_1509;
      ptr_deref_1521_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1521_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1521_root_address_inst_ack_0 <= ptr_deref_1521_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1521_resized_base_address;
      ptr_deref_1521_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1545_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1545_addr_0_ack_0 <= ptr_deref_1545_addr_0_req_0;
      aggregated_sig <= ptr_deref_1545_root_address;
      ptr_deref_1545_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1545_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1545_gather_scatter_ack_0 <= ptr_deref_1545_gather_scatter_req_0;
      aggregated_sig <= tmp63_1533;
      ptr_deref_1545_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1545_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1545_root_address_inst_ack_0 <= ptr_deref_1545_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1545_resized_base_address;
      ptr_deref_1545_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1569_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1569_addr_0_ack_0 <= ptr_deref_1569_addr_0_req_0;
      aggregated_sig <= ptr_deref_1569_root_address;
      ptr_deref_1569_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1569_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1569_gather_scatter_ack_0 <= ptr_deref_1569_gather_scatter_req_0;
      aggregated_sig <= tmp66_1557;
      ptr_deref_1569_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1569_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1569_root_address_inst_ack_0 <= ptr_deref_1569_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1569_resized_base_address;
      ptr_deref_1569_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1587_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1587_addr_0_ack_0 <= ptr_deref_1587_addr_0_req_0;
      aggregated_sig <= ptr_deref_1587_root_address;
      ptr_deref_1587_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1587_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1587_gather_scatter_ack_0 <= ptr_deref_1587_gather_scatter_req_0;
      aggregated_sig <= tmp68_1575;
      ptr_deref_1587_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1587_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1587_root_address_inst_ack_0 <= ptr_deref_1587_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1587_resized_base_address;
      ptr_deref_1587_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_969_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_969_gather_scatter_ack_0 <= ptr_deref_969_gather_scatter_req_0;
      aggregated_sig <= type_cast_971_wire_constant;
      ptr_deref_969_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    if_stmt_1000_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp2x_xi_999;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1000_branch_req_0,
          ack0 => if_stmt_1000_branch_ack_0,
          ack1 => if_stmt_1000_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1167_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1169_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1167_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_1167_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1167_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1172_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1167_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_1167_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1167_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_1169_wire_constant_cmp & expr_1172_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1167_branch_default_req_0,
          ack0 => switch_stmt_1167_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1028_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1028_resized_base_address;
      array_obj_ref_1028_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000001000",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1028_root_address_inst_req_0,
          ackL => array_obj_ref_1028_root_address_inst_ack_0,
          reqR => array_obj_ref_1028_root_address_inst_req_1,
          ackR => array_obj_ref_1028_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1102_root_address_inst array_obj_ref_1033_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1102_resized_base_address & array_obj_ref_1033_resized_base_address;
      array_obj_ref_1102_root_address <= data_out(21 downto 11);
      array_obj_ref_1033_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1102_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1033_root_address_inst_req_0;
      array_obj_ref_1102_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1033_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1102_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1033_root_address_inst_req_1;
      array_obj_ref_1102_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1033_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1038_root_address_inst array_obj_ref_1107_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1038_resized_base_address & array_obj_ref_1107_resized_base_address;
      array_obj_ref_1038_root_address <= data_out(21 downto 11);
      array_obj_ref_1107_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1038_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1107_root_address_inst_req_0;
      array_obj_ref_1038_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1107_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1038_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1107_root_address_inst_req_1;
      array_obj_ref_1038_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1107_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000010",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1043_root_address_inst array_obj_ref_1112_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1043_resized_base_address & array_obj_ref_1112_resized_base_address;
      array_obj_ref_1043_root_address <= data_out(21 downto 11);
      array_obj_ref_1112_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1043_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1112_root_address_inst_req_0;
      array_obj_ref_1043_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1112_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1043_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1112_root_address_inst_req_1;
      array_obj_ref_1043_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1112_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000011",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1048_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1048_resized_base_address;
      array_obj_ref_1048_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1048_root_address_inst_req_0,
          ackL => array_obj_ref_1048_root_address_inst_ack_0,
          reqR => array_obj_ref_1048_root_address_inst_req_1,
          ackR => array_obj_ref_1048_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1057_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1057_resized_base_address;
      array_obj_ref_1057_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000101",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1057_root_address_inst_req_0,
          ackL => array_obj_ref_1057_root_address_inst_ack_0,
          reqR => array_obj_ref_1057_root_address_inst_req_1,
          ackR => array_obj_ref_1057_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1062_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1062_resized_base_address;
      array_obj_ref_1062_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000110",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1062_root_address_inst_req_0,
          ackL => array_obj_ref_1062_root_address_inst_ack_0,
          reqR => array_obj_ref_1062_root_address_inst_req_1,
          ackR => array_obj_ref_1062_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_1067_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1067_resized_base_address;
      array_obj_ref_1067_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000111",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1067_root_address_inst_req_0,
          ackL => array_obj_ref_1067_root_address_inst_ack_0,
          reqR => array_obj_ref_1067_root_address_inst_req_1,
          ackR => array_obj_ref_1067_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_1093_index_0_scale 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1092_resized;
      simple_obj_ref_1092_scaled <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1093_index_0_scale_req_0,
          ackL => array_obj_ref_1093_index_0_scale_ack_0,
          reqR => array_obj_ref_1093_index_0_scale_req_1,
          ackR => array_obj_ref_1093_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_1093_root_address_inst array_obj_ref_1422_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1093_final_offset & array_obj_ref_1093_resized_base_address & array_obj_ref_1422_final_offset & array_obj_ref_1422_resized_base_address;
      array_obj_ref_1093_root_address <= data_out(21 downto 11);
      array_obj_ref_1422_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1093_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1422_root_address_inst_req_0;
      array_obj_ref_1093_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1422_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1093_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1422_root_address_inst_req_1;
      array_obj_ref_1093_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1422_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_1122_index_0_scale 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1121_resized;
      simple_obj_ref_1121_scaled <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1122_index_0_scale_req_0,
          ackL => array_obj_ref_1122_index_0_scale_ack_0,
          reqR => array_obj_ref_1122_index_0_scale_req_1,
          ackR => array_obj_ref_1122_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_1446_root_address_inst array_obj_ref_1122_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1446_final_offset & array_obj_ref_1446_resized_base_address & array_obj_ref_1122_final_offset & array_obj_ref_1122_resized_base_address;
      array_obj_ref_1446_root_address <= data_out(21 downto 11);
      array_obj_ref_1122_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1446_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1122_root_address_inst_req_0;
      array_obj_ref_1446_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1122_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1446_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1122_root_address_inst_req_1;
      array_obj_ref_1446_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1122_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_1131_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1131_resized_base_address;
      array_obj_ref_1131_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1131_root_address_inst_req_0,
          ackL => array_obj_ref_1131_root_address_inst_ack_0,
          reqR => array_obj_ref_1131_root_address_inst_req_1,
          ackR => array_obj_ref_1131_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_1136_root_address_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1136_resized_base_address;
      array_obj_ref_1136_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000010",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1136_root_address_inst_req_0,
          ackL => array_obj_ref_1136_root_address_inst_ack_0,
          reqR => array_obj_ref_1136_root_address_inst_req_1,
          ackR => array_obj_ref_1136_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_1141_root_address_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1141_resized_base_address;
      array_obj_ref_1141_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000011",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1141_root_address_inst_req_0,
          ackL => array_obj_ref_1141_root_address_inst_ack_0,
          reqR => array_obj_ref_1141_root_address_inst_req_1,
          ackR => array_obj_ref_1141_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : array_obj_ref_1470_root_address_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1470_final_offset & array_obj_ref_1470_resized_base_address;
      array_obj_ref_1470_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1470_root_address_inst_req_0,
          ackL => array_obj_ref_1470_root_address_inst_ack_0,
          reqR => array_obj_ref_1470_root_address_inst_req_1,
          ackR => array_obj_ref_1470_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : array_obj_ref_1494_root_address_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1494_final_offset & array_obj_ref_1494_resized_base_address;
      array_obj_ref_1494_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1494_root_address_inst_req_0,
          ackL => array_obj_ref_1494_root_address_inst_ack_0,
          reqR => array_obj_ref_1494_root_address_inst_req_1,
          ackR => array_obj_ref_1494_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : array_obj_ref_1518_root_address_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1518_final_offset & array_obj_ref_1518_resized_base_address;
      array_obj_ref_1518_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1518_root_address_inst_req_0,
          ackL => array_obj_ref_1518_root_address_inst_ack_0,
          reqR => array_obj_ref_1518_root_address_inst_req_1,
          ackR => array_obj_ref_1518_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : array_obj_ref_1542_root_address_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1542_final_offset & array_obj_ref_1542_resized_base_address;
      array_obj_ref_1542_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1542_root_address_inst_req_0,
          ackL => array_obj_ref_1542_root_address_inst_ack_0,
          reqR => array_obj_ref_1542_root_address_inst_req_1,
          ackR => array_obj_ref_1542_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : array_obj_ref_1566_root_address_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1566_final_offset & array_obj_ref_1566_resized_base_address;
      array_obj_ref_1566_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1566_root_address_inst_req_0,
          ackL => array_obj_ref_1566_root_address_inst_ack_0,
          reqR => array_obj_ref_1566_root_address_inst_req_1,
          ackR => array_obj_ref_1566_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : array_obj_ref_1584_root_address_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1584_final_offset & array_obj_ref_1584_resized_base_address;
      array_obj_ref_1584_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1584_root_address_inst_req_0,
          ackL => array_obj_ref_1584_root_address_inst_ack_0,
          reqR => array_obj_ref_1584_root_address_inst_req_1,
          ackR => array_obj_ref_1584_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1083_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_9_1071;
      tmp_1084 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1083_inst_req_0,
          ackL => binary_1083_inst_ack_0,
          reqR => binary_1083_inst_req_1,
          ackR => binary_1083_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1089_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1084;
      tmp138_1090 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1089_inst_req_0,
          ackL => binary_1089_inst_ack_0,
          reqR => binary_1089_inst_req_1,
          ackR => binary_1089_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1118_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1084;
      tmp146_1119 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1118_inst_req_0,
          ackL => binary_1118_inst_ack_0,
          reqR => binary_1118_inst_req_1,
          ackR => binary_1118_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1182_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp1_1183 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1182_inst_req_0,
          ackL => binary_1182_inst_ack_0,
          reqR => binary_1182_inst_req_1,
          ackR => binary_1182_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1196_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp4_1197 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1196_inst_req_0,
          ackL => binary_1196_inst_ack_0,
          reqR => binary_1196_inst_req_1,
          ackR => binary_1196_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1210_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp7_1211 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1210_inst_req_0,
          ackL => binary_1210_inst_ack_0,
          reqR => binary_1210_inst_req_1,
          ackR => binary_1210_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_1224_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp10_1225 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1224_inst_req_0,
          ackL => binary_1224_inst_ack_0,
          reqR => binary_1224_inst_req_1,
          ackR => binary_1224_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_1238_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp13_1239 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1238_inst_req_0,
          ackL => binary_1238_inst_ack_0,
          reqR => binary_1238_inst_req_1,
          ackR => binary_1238_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_1252_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp16_1253 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1252_inst_req_0,
          ackL => binary_1252_inst_ack_0,
          reqR => binary_1252_inst_req_1,
          ackR => binary_1252_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_1266_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp19_1267 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1266_inst_req_0,
          ackL => binary_1266_inst_ack_0,
          reqR => binary_1266_inst_req_1,
          ackR => binary_1266_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_1290_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp24_1291 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1290_inst_req_0,
          ackL => binary_1290_inst_ack_0,
          reqR => binary_1290_inst_req_1,
          ackR => binary_1290_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_1304_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp27_1305 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1304_inst_req_0,
          ackL => binary_1304_inst_ack_0,
          reqR => binary_1304_inst_req_1,
          ackR => binary_1304_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_1318_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp30_1319 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1318_inst_req_0,
          ackL => binary_1318_inst_ack_0,
          reqR => binary_1318_inst_req_1,
          ackR => binary_1318_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_1332_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp33_1333 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1332_inst_req_0,
          ackL => binary_1332_inst_ack_0,
          reqR => binary_1332_inst_req_1,
          ackR => binary_1332_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_1346_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp36_1347 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1346_inst_req_0,
          ackL => binary_1346_inst_ack_0,
          reqR => binary_1346_inst_req_1,
          ackR => binary_1346_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_1360_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp39_1361 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1360_inst_req_0,
          ackL => binary_1360_inst_ack_0,
          reqR => binary_1360_inst_req_1,
          ackR => binary_1360_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_1374_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp42_1375 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1374_inst_req_0,
          ackL => binary_1374_inst_ack_0,
          reqR => binary_1374_inst_req_1,
          ackR => binary_1374_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_1396_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_9_1071;
      tmp110_1397 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1396_inst_req_0,
          ackL => binary_1396_inst_ack_0,
          reqR => binary_1396_inst_req_1,
          ackR => binary_1396_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_1408_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp47_1409 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1408_inst_req_0,
          ackL => binary_1408_inst_ack_0,
          reqR => binary_1408_inst_req_1,
          ackR => binary_1408_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_1418_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_9_1071;
      tmp112_1419 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1418_inst_req_0,
          ackL => binary_1418_inst_ack_0,
          reqR => binary_1418_inst_req_1,
          ackR => binary_1418_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_1432_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp50_1433 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1432_inst_req_0,
          ackL => binary_1432_inst_ack_0,
          reqR => binary_1432_inst_req_1,
          ackR => binary_1432_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_1442_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp112_1419;
      tmp115_1443 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1442_inst_req_0,
          ackL => binary_1442_inst_ack_0,
          reqR => binary_1442_inst_req_1,
          ackR => binary_1442_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_1456_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp53_1457 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1456_inst_req_0,
          ackL => binary_1456_inst_ack_0,
          reqR => binary_1456_inst_req_1,
          ackR => binary_1456_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_1466_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp112_1419;
      tmp118_1467 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1466_inst_req_0,
          ackL => binary_1466_inst_ack_0,
          reqR => binary_1466_inst_req_1,
          ackR => binary_1466_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_1480_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp56_1481 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1480_inst_req_0,
          ackL => binary_1480_inst_ack_0,
          reqR => binary_1480_inst_req_1,
          ackR => binary_1480_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_1490_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp112_1419;
      tmp121_1491 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1490_inst_req_0,
          ackL => binary_1490_inst_ack_0,
          reqR => binary_1490_inst_req_1,
          ackR => binary_1490_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_1504_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp59_1505 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1504_inst_req_0,
          ackL => binary_1504_inst_ack_0,
          reqR => binary_1504_inst_req_1,
          ackR => binary_1504_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_1514_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp112_1419;
      tmp124_1515 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1514_inst_req_0,
          ackL => binary_1514_inst_ack_0,
          reqR => binary_1514_inst_req_1,
          ackR => binary_1514_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_1528_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp62_1529 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1528_inst_req_0,
          ackL => binary_1528_inst_ack_0,
          reqR => binary_1528_inst_req_1,
          ackR => binary_1528_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_1538_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp112_1419;
      tmp127_1539 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1538_inst_req_0,
          ackL => binary_1538_inst_ack_0,
          reqR => binary_1538_inst_req_1,
          ackR => binary_1538_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_1552_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1153;
      tmp65_1553 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1552_inst_req_0,
          ackL => binary_1552_inst_ack_0,
          reqR => binary_1552_inst_req_1,
          ackR => binary_1552_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_1562_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp112_1419;
      tmp130_1563 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1562_inst_req_0,
          ackL => binary_1562_inst_ack_0,
          reqR => binary_1562_inst_req_1,
          ackR => binary_1562_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : binary_1580_inst 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp112_1419;
      tmp133_1581 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1580_inst_req_0,
          ackL => binary_1580_inst_ack_0,
          reqR => binary_1580_inst_req_1,
          ackR => binary_1580_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : binary_998_inst 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xi_993;
      tmp2x_xi_999 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_998_inst_req_0,
          ackL => binary_998_inst_ack_0,
          reqR => binary_998_inst_req_1,
          ackR => binary_998_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : switch_stmt_1167_select_expr_0 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp76_1166;
      expr_1169_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_1167_select_expr_0_req_0,
          ackL => switch_stmt_1167_select_expr_0_ack_0,
          reqR => switch_stmt_1167_select_expr_0_req_1,
          ackR => switch_stmt_1167_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : switch_stmt_1167_select_expr_1 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp76_1166;
      expr_1172_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_1167_select_expr_1_req_0,
          ackL => switch_stmt_1167_select_expr_1_ack_0,
          reqR => switch_stmt_1167_select_expr_1_req_1,
          ackR => switch_stmt_1167_select_expr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared store operator group (0) : ptr_deref_1189_store_0 ptr_deref_1297_store_0 ptr_deref_1425_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1189_store_0_req_0;
      reqL(1) <= ptr_deref_1297_store_0_req_0;
      reqL(0) <= ptr_deref_1425_store_0_req_0;
      ptr_deref_1189_store_0_ack_0 <= ackL(2);
      ptr_deref_1297_store_0_ack_0 <= ackL(1);
      ptr_deref_1425_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1189_store_0_req_1;
      reqR(1) <= ptr_deref_1297_store_0_req_1;
      reqR(0) <= ptr_deref_1425_store_0_req_1;
      ptr_deref_1189_store_0_ack_1 <= ackR(2);
      ptr_deref_1297_store_0_ack_1 <= ackR(1);
      ptr_deref_1425_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1189_word_address_0 & ptr_deref_1297_word_address_0 & ptr_deref_1425_word_address_0;
      data_in <= ptr_deref_1189_data_0 & ptr_deref_1297_data_0 & ptr_deref_1425_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(7),
          mack => memory_space_0_sr_ack(7),
          maddr => memory_space_0_sr_addr(87 downto 77),
          mdata => memory_space_0_sr_data(63 downto 56),
          mtag => memory_space_0_sr_tag(15 downto 14),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(7),
          mack => memory_space_0_sc_ack(7),
          mtag => memory_space_0_sc_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1203_store_0 ptr_deref_1311_store_0 ptr_deref_1449_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1203_store_0_req_0;
      reqL(1) <= ptr_deref_1311_store_0_req_0;
      reqL(0) <= ptr_deref_1449_store_0_req_0;
      ptr_deref_1203_store_0_ack_0 <= ackL(2);
      ptr_deref_1311_store_0_ack_0 <= ackL(1);
      ptr_deref_1449_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1203_store_0_req_1;
      reqR(1) <= ptr_deref_1311_store_0_req_1;
      reqR(0) <= ptr_deref_1449_store_0_req_1;
      ptr_deref_1203_store_0_ack_1 <= ackR(2);
      ptr_deref_1311_store_0_ack_1 <= ackR(1);
      ptr_deref_1449_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1203_word_address_0 & ptr_deref_1311_word_address_0 & ptr_deref_1449_word_address_0;
      data_in <= ptr_deref_1203_data_0 & ptr_deref_1311_data_0 & ptr_deref_1449_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(6),
          mack => memory_space_0_sr_ack(6),
          maddr => memory_space_0_sr_addr(76 downto 66),
          mdata => memory_space_0_sr_data(55 downto 48),
          mtag => memory_space_0_sr_tag(13 downto 12),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(6),
          mack => memory_space_0_sc_ack(6),
          mtag => memory_space_0_sc_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_1217_store_0 ptr_deref_1325_store_0 ptr_deref_1473_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1217_store_0_req_0;
      reqL(1) <= ptr_deref_1325_store_0_req_0;
      reqL(0) <= ptr_deref_1473_store_0_req_0;
      ptr_deref_1217_store_0_ack_0 <= ackL(2);
      ptr_deref_1325_store_0_ack_0 <= ackL(1);
      ptr_deref_1473_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1217_store_0_req_1;
      reqR(1) <= ptr_deref_1325_store_0_req_1;
      reqR(0) <= ptr_deref_1473_store_0_req_1;
      ptr_deref_1217_store_0_ack_1 <= ackR(2);
      ptr_deref_1325_store_0_ack_1 <= ackR(1);
      ptr_deref_1473_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1217_word_address_0 & ptr_deref_1325_word_address_0 & ptr_deref_1473_word_address_0;
      data_in <= ptr_deref_1217_data_0 & ptr_deref_1325_data_0 & ptr_deref_1473_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(5),
          mack => memory_space_0_sr_ack(5),
          maddr => memory_space_0_sr_addr(65 downto 55),
          mdata => memory_space_0_sr_data(47 downto 40),
          mtag => memory_space_0_sr_tag(11 downto 10),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(5),
          mack => memory_space_0_sc_ack(5),
          mtag => memory_space_0_sc_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_1339_store_0 ptr_deref_1231_store_0 ptr_deref_1497_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1339_store_0_req_0;
      reqL(1) <= ptr_deref_1231_store_0_req_0;
      reqL(0) <= ptr_deref_1497_store_0_req_0;
      ptr_deref_1339_store_0_ack_0 <= ackL(2);
      ptr_deref_1231_store_0_ack_0 <= ackL(1);
      ptr_deref_1497_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1339_store_0_req_1;
      reqR(1) <= ptr_deref_1231_store_0_req_1;
      reqR(0) <= ptr_deref_1497_store_0_req_1;
      ptr_deref_1339_store_0_ack_1 <= ackR(2);
      ptr_deref_1231_store_0_ack_1 <= ackR(1);
      ptr_deref_1497_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1339_word_address_0 & ptr_deref_1231_word_address_0 & ptr_deref_1497_word_address_0;
      data_in <= ptr_deref_1339_data_0 & ptr_deref_1231_data_0 & ptr_deref_1497_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(4),
          mack => memory_space_0_sr_ack(4),
          maddr => memory_space_0_sr_addr(54 downto 44),
          mdata => memory_space_0_sr_data(39 downto 32),
          mtag => memory_space_0_sr_tag(9 downto 8),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(4),
          mack => memory_space_0_sc_ack(4),
          mtag => memory_space_0_sc_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_1245_store_0 ptr_deref_1353_store_0 ptr_deref_1521_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1245_store_0_req_0;
      reqL(1) <= ptr_deref_1353_store_0_req_0;
      reqL(0) <= ptr_deref_1521_store_0_req_0;
      ptr_deref_1245_store_0_ack_0 <= ackL(2);
      ptr_deref_1353_store_0_ack_0 <= ackL(1);
      ptr_deref_1521_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1245_store_0_req_1;
      reqR(1) <= ptr_deref_1353_store_0_req_1;
      reqR(0) <= ptr_deref_1521_store_0_req_1;
      ptr_deref_1245_store_0_ack_1 <= ackR(2);
      ptr_deref_1353_store_0_ack_1 <= ackR(1);
      ptr_deref_1521_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1245_word_address_0 & ptr_deref_1353_word_address_0 & ptr_deref_1521_word_address_0;
      data_in <= ptr_deref_1245_data_0 & ptr_deref_1353_data_0 & ptr_deref_1521_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(3),
          mack => memory_space_0_sr_ack(3),
          maddr => memory_space_0_sr_addr(43 downto 33),
          mdata => memory_space_0_sr_data(31 downto 24),
          mtag => memory_space_0_sr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(3),
          mack => memory_space_0_sc_ack(3),
          mtag => memory_space_0_sc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_1367_store_0 ptr_deref_1259_store_0 ptr_deref_1545_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1367_store_0_req_0;
      reqL(1) <= ptr_deref_1259_store_0_req_0;
      reqL(0) <= ptr_deref_1545_store_0_req_0;
      ptr_deref_1367_store_0_ack_0 <= ackL(2);
      ptr_deref_1259_store_0_ack_0 <= ackL(1);
      ptr_deref_1545_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1367_store_0_req_1;
      reqR(1) <= ptr_deref_1259_store_0_req_1;
      reqR(0) <= ptr_deref_1545_store_0_req_1;
      ptr_deref_1367_store_0_ack_1 <= ackR(2);
      ptr_deref_1259_store_0_ack_1 <= ackR(1);
      ptr_deref_1545_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1367_word_address_0 & ptr_deref_1259_word_address_0 & ptr_deref_1545_word_address_0;
      data_in <= ptr_deref_1367_data_0 & ptr_deref_1259_data_0 & ptr_deref_1545_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(2),
          mack => memory_space_0_sr_ack(2),
          maddr => memory_space_0_sr_addr(32 downto 22),
          mdata => memory_space_0_sr_data(23 downto 16),
          mtag => memory_space_0_sr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(2),
          mack => memory_space_0_sc_ack(2),
          mtag => memory_space_0_sc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_1381_store_0 ptr_deref_1273_store_0 ptr_deref_1569_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1381_store_0_req_0;
      reqL(1) <= ptr_deref_1273_store_0_req_0;
      reqL(0) <= ptr_deref_1569_store_0_req_0;
      ptr_deref_1381_store_0_ack_0 <= ackL(2);
      ptr_deref_1273_store_0_ack_0 <= ackL(1);
      ptr_deref_1569_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1381_store_0_req_1;
      reqR(1) <= ptr_deref_1273_store_0_req_1;
      reqR(0) <= ptr_deref_1569_store_0_req_1;
      ptr_deref_1381_store_0_ack_1 <= ackR(2);
      ptr_deref_1273_store_0_ack_1 <= ackR(1);
      ptr_deref_1569_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1381_word_address_0 & ptr_deref_1273_word_address_0 & ptr_deref_1569_word_address_0;
      data_in <= ptr_deref_1381_data_0 & ptr_deref_1273_data_0 & ptr_deref_1569_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(1),
          mack => memory_space_0_sr_ack(1),
          maddr => memory_space_0_sr_addr(21 downto 11),
          mdata => memory_space_0_sr_data(15 downto 8),
          mtag => memory_space_0_sr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(1),
          mack => memory_space_0_sc_ack(1),
          mtag => memory_space_0_sc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_1281_store_0 ptr_deref_1389_store_0 ptr_deref_1587_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1281_store_0_req_0;
      reqL(1) <= ptr_deref_1389_store_0_req_0;
      reqL(0) <= ptr_deref_1587_store_0_req_0;
      ptr_deref_1281_store_0_ack_0 <= ackL(2);
      ptr_deref_1389_store_0_ack_0 <= ackL(1);
      ptr_deref_1587_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1281_store_0_req_1;
      reqR(1) <= ptr_deref_1389_store_0_req_1;
      reqR(0) <= ptr_deref_1587_store_0_req_1;
      ptr_deref_1281_store_0_ack_1 <= ackR(2);
      ptr_deref_1389_store_0_ack_1 <= ackR(1);
      ptr_deref_1587_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1281_word_address_0 & ptr_deref_1389_word_address_0 & ptr_deref_1587_word_address_0;
      data_in <= ptr_deref_1281_data_0 & ptr_deref_1389_data_0 & ptr_deref_1587_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(10 downto 0),
          mdata => memory_space_0_sr_data(7 downto 0),
          mtag => memory_space_0_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared store operator group (8) : ptr_deref_969_store_0 
    StoreGroup8: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_969_store_0_req_0;
      ptr_deref_969_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_969_store_0_req_1;
      ptr_deref_969_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_969_word_address_0;
      data_in <= ptr_deref_969_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(3 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 8
    -- shared inport operator group (0) : simple_obj_ref_1014_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1014_inst_req_0;
      simple_obj_ref_1014_inst_ack_0 <= ack(0);
      tmp4x_xi_1015 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_get_pipe_read_req(0),
          oack => free_queue_get_pipe_read_ack(0),
          odata => free_queue_get_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_1152_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1152_inst_req_0;
      simple_obj_ref_1152_inst_ack_0 <= ack(0);
      tmp74_1153 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_1161_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1161_inst_req_0;
      simple_obj_ref_1161_inst_ack_0 <= ack(0);
      tmp75_1162 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_ctrl_pipe_read_req(0),
          oack => in_ctrl_pipe_read_ack(0),
          odata => in_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_992_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_992_inst_req_0;
      simple_obj_ref_992_inst_ack_0 <= ack(0);
      tmpx_xi_993 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_ack_pipe_read_req(0),
          oack => free_queue_ack_pipe_read_ack(0),
          odata => free_queue_ack_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : simple_obj_ref_1596_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1596_inst_req_0;
      simple_obj_ref_1596_inst_ack_0 <= ack(0);
      data_in <= tmp4x_xi_1015;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => midpipe_pipe_write_req(0),
          oack => midpipe_pipe_write_ack(0),
          odata => midpipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_981_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_981_inst_req_0;
      simple_obj_ref_981_inst_ack_0 <= ack(0);
      data_in <= type_cast_983_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_output is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_0_lr_req : out  std_logic_vector(7 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(7 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(87 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(15 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(7 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(7 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(15 downto 0);
    midpipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    midpipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    midpipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
    out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_output;
architecture Default of wrapper_output is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_output_CP_7359_start: Boolean;
  -- links between control-path and data-path
  signal binary_1783_inst_ack_0 : boolean;
  signal array_obj_ref_1858_index_0_resize_ack_0 : boolean;
  signal binary_1834_inst_ack_1 : boolean;
  signal binary_1793_inst_ack_0 : boolean;
  signal ptr_deref_1748_addr_0_req_0 : boolean;
  signal array_obj_ref_1848_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1748_addr_0_ack_0 : boolean;
  signal binary_1793_inst_req_0 : boolean;
  signal binary_1793_inst_ack_1 : boolean;
  signal ptr_deref_1748_load_0_ack_0 : boolean;
  signal ptr_deref_1639_load_0_ack_1 : boolean;
  signal simple_obj_ref_1811_inst_ack_0 : boolean;
  signal binary_1793_inst_req_1 : boolean;
  signal array_obj_ref_1838_index_0_resize_req_0 : boolean;
  signal binary_1783_inst_req_1 : boolean;
  signal ptr_deref_1639_base_resize_req_0 : boolean;
  signal binary_1788_inst_ack_1 : boolean;
  signal binary_1783_inst_ack_1 : boolean;
  signal ptr_deref_1748_root_address_inst_ack_0 : boolean;
  signal binary_1783_inst_req_0 : boolean;
  signal ptr_deref_1748_load_0_req_0 : boolean;
  signal array_obj_ref_1858_index_0_rename_req_0 : boolean;
  signal binary_1834_inst_req_1 : boolean;
  signal binary_1844_inst_ack_1 : boolean;
  signal simple_obj_ref_1801_inst_ack_0 : boolean;
  signal array_obj_ref_1848_base_resize_req_0 : boolean;
  signal ptr_deref_1748_root_address_inst_req_0 : boolean;
  signal binary_1763_inst_ack_1 : boolean;
  signal binary_1834_inst_ack_0 : boolean;
  signal binary_1844_inst_req_1 : boolean;
  signal binary_1763_inst_req_1 : boolean;
  signal binary_1768_inst_ack_1 : boolean;
  signal ptr_deref_1748_load_0_ack_1 : boolean;
  signal binary_1864_inst_req_1 : boolean;
  signal ptr_deref_1748_gather_scatter_ack_0 : boolean;
  signal binary_1844_inst_ack_0 : boolean;
  signal binary_1768_inst_ack_0 : boolean;
  signal ptr_deref_1639_base_resize_ack_0 : boolean;
  signal binary_1768_inst_req_1 : boolean;
  signal simple_obj_ref_1801_inst_req_0 : boolean;
  signal binary_2019_inst_ack_0 : boolean;
  signal ptr_deref_1639_gather_scatter_ack_0 : boolean;
  signal binary_1763_inst_ack_0 : boolean;
  signal binary_1844_inst_req_0 : boolean;
  signal binary_1763_inst_req_0 : boolean;
  signal binary_1788_inst_req_1 : boolean;
  signal binary_1788_inst_ack_0 : boolean;
  signal array_obj_ref_1654_final_reg_req_0 : boolean;
  signal array_obj_ref_1635_final_reg_ack_0 : boolean;
  signal array_obj_ref_1858_base_resize_req_0 : boolean;
  signal binary_1834_inst_req_0 : boolean;
  signal ptr_deref_1748_base_resize_req_0 : boolean;
  signal array_obj_ref_1848_root_address_inst_req_1 : boolean;
  signal binary_1788_inst_req_0 : boolean;
  signal array_obj_ref_1858_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1748_base_resize_ack_0 : boolean;
  signal binary_1778_inst_req_1 : boolean;
  signal ptr_deref_1639_root_address_inst_req_0 : boolean;
  signal ptr_deref_1748_gather_scatter_req_0 : boolean;
  signal ptr_deref_1639_addr_0_ack_0 : boolean;
  signal binary_1668_inst_req_1 : boolean;
  signal array_obj_ref_1744_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1848_offset_inst_req_0 : boolean;
  signal ptr_deref_1658_root_address_inst_req_0 : boolean;
  signal binary_1768_inst_req_0 : boolean;
  signal array_obj_ref_1838_final_reg_ack_0 : boolean;
  signal ptr_deref_1934_addr_0_req_0 : boolean;
  signal binary_1778_inst_ack_0 : boolean;
  signal array_obj_ref_1654_final_reg_ack_0 : boolean;
  signal array_obj_ref_1673_root_address_inst_ack_1 : boolean;
  signal binary_1864_inst_req_0 : boolean;
  signal array_obj_ref_1858_index_0_resize_req_0 : boolean;
  signal ptr_deref_1658_addr_0_req_0 : boolean;
  signal ptr_deref_1639_load_0_req_1 : boolean;
  signal array_obj_ref_1744_final_reg_ack_0 : boolean;
  signal array_obj_ref_1848_base_resize_ack_0 : boolean;
  signal binary_1758_inst_ack_1 : boolean;
  signal type_cast_1630_inst_req_0 : boolean;
  signal array_obj_ref_1858_base_resize_ack_0 : boolean;
  signal type_cast_1643_inst_ack_0 : boolean;
  signal ptr_deref_1658_gather_scatter_req_0 : boolean;
  signal ptr_deref_1658_base_resize_req_0 : boolean;
  signal binary_1668_inst_ack_1 : boolean;
  signal binary_1758_inst_req_1 : boolean;
  signal binary_1854_inst_req_1 : boolean;
  signal array_obj_ref_1858_final_reg_req_0 : boolean;
  signal type_cast_1643_inst_req_0 : boolean;
  signal type_cast_1630_inst_ack_0 : boolean;
  signal ptr_deref_1658_addr_0_ack_0 : boolean;
  signal type_cast_1662_inst_req_0 : boolean;
  signal array_obj_ref_1744_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1639_addr_0_req_0 : boolean;
  signal array_obj_ref_1635_base_resize_req_0 : boolean;
  signal ptr_deref_1658_load_0_req_1 : boolean;
  signal array_obj_ref_1635_base_resize_ack_0 : boolean;
  signal ptr_deref_1639_load_0_req_0 : boolean;
  signal array_obj_ref_1858_final_reg_ack_0 : boolean;
  signal type_cast_1662_inst_ack_0 : boolean;
  signal binary_1758_inst_req_0 : boolean;
  signal binary_1778_inst_ack_1 : boolean;
  signal ptr_deref_1639_load_0_ack_0 : boolean;
  signal binary_1778_inst_req_0 : boolean;
  signal array_obj_ref_1635_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1838_final_reg_req_0 : boolean;
  signal ptr_deref_1658_load_0_ack_1 : boolean;
  signal array_obj_ref_1838_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1838_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1848_offset_inst_ack_0 : boolean;
  signal binary_1854_inst_req_0 : boolean;
  signal binary_1854_inst_ack_1 : boolean;
  signal binary_1758_inst_ack_0 : boolean;
  signal ptr_deref_1658_load_0_req_0 : boolean;
  signal array_obj_ref_1848_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1658_load_0_ack_0 : boolean;
  signal array_obj_ref_1868_index_0_resize_req_0 : boolean;
  signal ptr_deref_1639_root_address_inst_ack_0 : boolean;
  signal binary_1649_inst_req_0 : boolean;
  signal ptr_deref_1658_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1838_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1858_root_address_inst_req_1 : boolean;
  signal binary_1668_inst_req_0 : boolean;
  signal binary_1649_inst_ack_0 : boolean;
  signal ptr_deref_1677_load_0_req_0 : boolean;
  signal ptr_deref_1677_load_0_ack_0 : boolean;
  signal binary_1649_inst_req_1 : boolean;
  signal ptr_deref_1658_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1673_base_resize_req_0 : boolean;
  signal binary_1828_inst_ack_1 : boolean;
  signal binary_1649_inst_ack_1 : boolean;
  signal array_obj_ref_1838_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1673_base_resize_ack_0 : boolean;
  signal binary_1773_inst_req_0 : boolean;
  signal array_obj_ref_1848_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1848_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1838_index_0_rename_req_0 : boolean;
  signal ptr_deref_1677_addr_0_req_0 : boolean;
  signal array_obj_ref_1635_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1654_root_address_inst_req_0 : boolean;
  signal ptr_deref_1658_base_resize_ack_0 : boolean;
  signal array_obj_ref_1654_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1654_base_resize_req_0 : boolean;
  signal binary_2024_inst_ack_0 : boolean;
  signal array_obj_ref_1848_index_0_resize_ack_0 : boolean;
  signal type_cast_1752_inst_ack_0 : boolean;
  signal array_obj_ref_1858_root_address_inst_req_0 : boolean;
  signal ptr_deref_1639_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1838_offset_inst_req_0 : boolean;
  signal ptr_deref_1677_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1635_root_address_inst_req_1 : boolean;
  signal binary_1854_inst_ack_0 : boolean;
  signal array_obj_ref_1858_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1654_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1838_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1677_root_address_inst_req_0 : boolean;
  signal ptr_deref_1677_base_resize_req_0 : boolean;
  signal binary_1828_inst_req_0 : boolean;
  signal ptr_deref_1677_base_resize_ack_0 : boolean;
  signal array_obj_ref_1868_index_0_resize_ack_0 : boolean;
  signal binary_1828_inst_ack_0 : boolean;
  signal binary_1864_inst_ack_1 : boolean;
  signal ptr_deref_1677_addr_0_ack_0 : boolean;
  signal array_obj_ref_1848_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1635_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1673_root_address_inst_req_0 : boolean;
  signal binary_1828_inst_req_1 : boolean;
  signal array_obj_ref_1654_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1673_root_address_inst_ack_0 : boolean;
  signal binary_1773_inst_ack_1 : boolean;
  signal array_obj_ref_1838_base_resize_ack_0 : boolean;
  signal binary_1773_inst_req_1 : boolean;
  signal array_obj_ref_1673_final_reg_req_0 : boolean;
  signal array_obj_ref_1673_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1744_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1838_base_resize_req_0 : boolean;
  signal array_obj_ref_1654_base_resize_ack_0 : boolean;
  signal binary_1668_inst_ack_0 : boolean;
  signal array_obj_ref_1744_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1838_offset_inst_ack_0 : boolean;
  signal binary_1773_inst_ack_0 : boolean;
  signal array_obj_ref_1673_final_reg_ack_0 : boolean;
  signal array_obj_ref_1848_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1744_final_reg_req_0 : boolean;
  signal array_obj_ref_1635_final_reg_req_0 : boolean;
  signal ptr_deref_1934_root_address_inst_req_0 : boolean;
  signal ptr_deref_1677_load_0_req_1 : boolean;
  signal array_obj_ref_1838_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1677_load_0_ack_1 : boolean;
  signal ptr_deref_1677_gather_scatter_req_0 : boolean;
  signal ptr_deref_1677_gather_scatter_ack_0 : boolean;
  signal binary_2029_inst_ack_1 : boolean;
  signal array_obj_ref_1858_offset_inst_req_0 : boolean;
  signal array_obj_ref_1858_offset_inst_ack_0 : boolean;
  signal ptr_deref_1976_addr_0_ack_0 : boolean;
  signal ptr_deref_1976_addr_0_req_0 : boolean;
  signal if_stmt_2063_branch_req_0 : boolean;
  signal array_obj_ref_1878_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1878_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1948_load_0_ack_0 : boolean;
  signal array_obj_ref_1878_index_0_rename_req_0 : boolean;
  signal binary_2014_inst_ack_1 : boolean;
  signal array_obj_ref_1878_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1948_load_0_req_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1948_load_0_ack_1 : boolean;
  signal ptr_deref_1990_base_resize_req_0 : boolean;
  signal array_obj_ref_1868_base_resize_ack_0 : boolean;
  signal binary_2019_inst_req_1 : boolean;
  signal ptr_deref_1976_load_0_ack_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_req_1 : boolean;
  signal binary_2024_inst_ack_1 : boolean;
  signal ptr_deref_1934_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1868_index_0_rename_req_0 : boolean;
  signal ptr_deref_1948_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_req_0 : boolean;
  signal binary_1864_inst_ack_0 : boolean;
  signal array_obj_ref_1868_base_resize_req_0 : boolean;
  signal array_obj_ref_1868_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1868_offset_inst_req_0 : boolean;
  signal ptr_deref_1948_load_0_req_1 : boolean;
  signal ptr_deref_1976_root_address_inst_req_0 : boolean;
  signal binary_2039_inst_ack_1 : boolean;
  signal array_obj_ref_1858_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1868_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1848_final_reg_req_0 : boolean;
  signal binary_2024_inst_req_0 : boolean;
  signal array_obj_ref_1848_final_reg_ack_0 : boolean;
  signal binary_1874_inst_req_1 : boolean;
  signal ptr_deref_1934_base_resize_ack_0 : boolean;
  signal binary_1874_inst_ack_1 : boolean;
  signal type_cast_1752_inst_req_0 : boolean;
  signal simple_obj_ref_1811_inst_req_0 : boolean;
  signal array_obj_ref_1868_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1868_final_reg_req_0 : boolean;
  signal ptr_deref_1976_load_0_req_0 : boolean;
  signal array_obj_ref_1868_final_reg_ack_0 : boolean;
  signal binary_1874_inst_req_0 : boolean;
  signal binary_1874_inst_ack_0 : boolean;
  signal ptr_deref_1748_load_0_req_1 : boolean;
  signal simple_obj_ref_1613_inst_req_0 : boolean;
  signal simple_obj_ref_1613_inst_ack_0 : boolean;
  signal type_cast_1617_inst_req_0 : boolean;
  signal type_cast_1617_inst_ack_0 : boolean;
  signal array_obj_ref_1622_base_resize_req_0 : boolean;
  signal array_obj_ref_1622_base_resize_ack_0 : boolean;
  signal array_obj_ref_1622_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1622_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1622_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1622_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1622_final_reg_req_0 : boolean;
  signal array_obj_ref_1622_final_reg_ack_0 : boolean;
  signal ptr_deref_1626_base_resize_req_0 : boolean;
  signal ptr_deref_1626_base_resize_ack_0 : boolean;
  signal ptr_deref_1626_root_address_inst_req_0 : boolean;
  signal ptr_deref_1626_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1626_addr_0_req_0 : boolean;
  signal ptr_deref_1626_addr_0_ack_0 : boolean;
  signal ptr_deref_1626_load_0_req_0 : boolean;
  signal ptr_deref_1626_load_0_ack_0 : boolean;
  signal ptr_deref_1626_load_0_req_1 : boolean;
  signal ptr_deref_1626_load_0_ack_1 : boolean;
  signal ptr_deref_1626_gather_scatter_req_0 : boolean;
  signal ptr_deref_1626_gather_scatter_ack_0 : boolean;
  signal binary_2024_inst_req_1 : boolean;
  signal type_cast_1681_inst_req_0 : boolean;
  signal type_cast_1681_inst_ack_0 : boolean;
  signal binary_2019_inst_ack_1 : boolean;
  signal binary_1958_inst_req_0 : boolean;
  signal binary_1687_inst_req_0 : boolean;
  signal binary_1687_inst_ack_0 : boolean;
  signal ptr_deref_1934_addr_0_ack_0 : boolean;
  signal binary_1687_inst_req_1 : boolean;
  signal binary_1687_inst_ack_1 : boolean;
  signal binary_2039_inst_req_0 : boolean;
  signal binary_2039_inst_ack_0 : boolean;
  signal ptr_deref_1948_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1692_base_resize_req_0 : boolean;
  signal array_obj_ref_1692_base_resize_ack_0 : boolean;
  signal binary_2029_inst_req_0 : boolean;
  signal array_obj_ref_1692_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1692_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1692_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1692_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1692_final_reg_req_0 : boolean;
  signal array_obj_ref_1692_final_reg_ack_0 : boolean;
  signal ptr_deref_1976_load_0_req_1 : boolean;
  signal ptr_deref_1696_base_resize_req_0 : boolean;
  signal ptr_deref_1976_load_0_ack_1 : boolean;
  signal ptr_deref_1696_base_resize_ack_0 : boolean;
  signal ptr_deref_1990_base_resize_ack_0 : boolean;
  signal ptr_deref_1696_root_address_inst_req_0 : boolean;
  signal ptr_deref_1976_gather_scatter_req_0 : boolean;
  signal ptr_deref_1696_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1696_addr_0_req_0 : boolean;
  signal ptr_deref_1696_addr_0_ack_0 : boolean;
  signal binary_2029_inst_ack_0 : boolean;
  signal ptr_deref_1696_load_0_req_0 : boolean;
  signal ptr_deref_1696_load_0_ack_0 : boolean;
  signal ptr_deref_1976_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1696_load_0_req_1 : boolean;
  signal ptr_deref_1696_load_0_ack_1 : boolean;
  signal ptr_deref_1696_gather_scatter_req_0 : boolean;
  signal ptr_deref_1696_gather_scatter_ack_0 : boolean;
  signal binary_2039_inst_req_1 : boolean;
  signal binary_2029_inst_req_1 : boolean;
  signal type_cast_1700_inst_req_0 : boolean;
  signal type_cast_1700_inst_ack_0 : boolean;
  signal binary_1706_inst_req_0 : boolean;
  signal binary_1706_inst_ack_0 : boolean;
  signal binary_1706_inst_req_1 : boolean;
  signal binary_1706_inst_ack_1 : boolean;
  signal type_cast_1980_inst_req_0 : boolean;
  signal type_cast_1952_inst_req_0 : boolean;
  signal type_cast_1980_inst_ack_0 : boolean;
  signal array_obj_ref_1711_base_resize_req_0 : boolean;
  signal array_obj_ref_1711_base_resize_ack_0 : boolean;
  signal array_obj_ref_1711_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1711_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1934_load_0_req_0 : boolean;
  signal array_obj_ref_1711_root_address_inst_req_1 : boolean;
  signal ptr_deref_1934_load_0_ack_0 : boolean;
  signal array_obj_ref_1711_root_address_inst_ack_1 : boolean;
  signal binary_1958_inst_ack_0 : boolean;
  signal array_obj_ref_1711_final_reg_req_0 : boolean;
  signal array_obj_ref_1711_final_reg_ack_0 : boolean;
  signal type_cast_1952_inst_ack_0 : boolean;
  signal binary_1986_inst_req_0 : boolean;
  signal binary_1986_inst_ack_0 : boolean;
  signal binary_1986_inst_req_1 : boolean;
  signal binary_1986_inst_ack_1 : boolean;
  signal ptr_deref_1715_base_resize_req_0 : boolean;
  signal ptr_deref_1990_root_address_inst_req_0 : boolean;
  signal binary_2019_inst_req_0 : boolean;
  signal ptr_deref_1715_base_resize_ack_0 : boolean;
  signal ptr_deref_1715_root_address_inst_req_0 : boolean;
  signal ptr_deref_1990_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1715_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1715_addr_0_req_0 : boolean;
  signal ptr_deref_1715_addr_0_ack_0 : boolean;
  signal ptr_deref_1715_load_0_req_0 : boolean;
  signal ptr_deref_1715_load_0_ack_0 : boolean;
  signal ptr_deref_1715_load_0_req_1 : boolean;
  signal ptr_deref_1715_load_0_ack_1 : boolean;
  signal ptr_deref_1715_gather_scatter_req_0 : boolean;
  signal ptr_deref_1715_gather_scatter_ack_0 : boolean;
  signal type_cast_1719_inst_req_0 : boolean;
  signal type_cast_1719_inst_ack_0 : boolean;
  signal binary_1725_inst_req_0 : boolean;
  signal binary_1725_inst_ack_0 : boolean;
  signal binary_1725_inst_req_1 : boolean;
  signal binary_1725_inst_ack_1 : boolean;
  signal ptr_deref_1729_base_resize_req_0 : boolean;
  signal ptr_deref_1729_base_resize_ack_0 : boolean;
  signal ptr_deref_1729_root_address_inst_req_0 : boolean;
  signal ptr_deref_1729_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1729_addr_0_req_0 : boolean;
  signal ptr_deref_1729_addr_0_ack_0 : boolean;
  signal ptr_deref_1729_load_0_req_0 : boolean;
  signal ptr_deref_1729_load_0_ack_0 : boolean;
  signal ptr_deref_1729_load_0_req_1 : boolean;
  signal ptr_deref_1729_load_0_ack_1 : boolean;
  signal ptr_deref_1729_gather_scatter_req_0 : boolean;
  signal ptr_deref_1729_gather_scatter_ack_0 : boolean;
  signal type_cast_1733_inst_req_0 : boolean;
  signal type_cast_1733_inst_ack_0 : boolean;
  signal binary_1739_inst_req_0 : boolean;
  signal binary_1739_inst_ack_0 : boolean;
  signal binary_1739_inst_req_1 : boolean;
  signal binary_1739_inst_ack_1 : boolean;
  signal array_obj_ref_1744_base_resize_req_0 : boolean;
  signal array_obj_ref_1744_base_resize_ack_0 : boolean;
  signal array_obj_ref_1878_offset_inst_req_0 : boolean;
  signal array_obj_ref_1878_offset_inst_ack_0 : boolean;
  signal ptr_deref_1976_root_address_inst_ack_0 : boolean;
  signal binary_2014_inst_req_1 : boolean;
  signal array_obj_ref_1878_base_resize_req_0 : boolean;
  signal array_obj_ref_1878_base_resize_ack_0 : boolean;
  signal binary_2014_inst_ack_0 : boolean;
  signal array_obj_ref_1878_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1878_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1878_root_address_inst_req_1 : boolean;
  signal ptr_deref_1934_base_resize_req_0 : boolean;
  signal binary_2014_inst_req_0 : boolean;
  signal array_obj_ref_1878_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1878_final_reg_req_0 : boolean;
  signal array_obj_ref_1878_final_reg_ack_0 : boolean;
  signal binary_2087_inst_req_0 : boolean;
  signal ptr_deref_1976_base_resize_ack_0 : boolean;
  signal ptr_deref_1976_base_resize_req_0 : boolean;
  signal ptr_deref_1948_addr_0_ack_0 : boolean;
  signal binary_1884_inst_req_0 : boolean;
  signal binary_1884_inst_ack_0 : boolean;
  signal binary_1884_inst_req_1 : boolean;
  signal binary_1884_inst_ack_1 : boolean;
  signal ptr_deref_1948_addr_0_req_0 : boolean;
  signal array_obj_ref_1888_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1888_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1948_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1888_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1888_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1948_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1888_offset_inst_req_0 : boolean;
  signal array_obj_ref_1888_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1888_base_resize_req_0 : boolean;
  signal array_obj_ref_1888_base_resize_ack_0 : boolean;
  signal binary_2087_inst_ack_1 : boolean;
  signal binary_1972_inst_ack_1 : boolean;
  signal array_obj_ref_1888_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1888_root_address_inst_ack_0 : boolean;
  signal binary_1972_inst_req_1 : boolean;
  signal array_obj_ref_1888_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1888_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1948_base_resize_ack_0 : boolean;
  signal array_obj_ref_1888_final_reg_req_0 : boolean;
  signal array_obj_ref_1888_final_reg_ack_0 : boolean;
  signal ptr_deref_1948_base_resize_req_0 : boolean;
  signal binary_1972_inst_ack_0 : boolean;
  signal binary_1972_inst_req_0 : boolean;
  signal binary_1894_inst_req_0 : boolean;
  signal binary_1894_inst_ack_0 : boolean;
  signal type_cast_2008_inst_ack_0 : boolean;
  signal binary_1894_inst_req_1 : boolean;
  signal type_cast_2008_inst_req_0 : boolean;
  signal binary_1894_inst_ack_1 : boolean;
  signal type_cast_1966_inst_ack_0 : boolean;
  signal type_cast_1966_inst_req_0 : boolean;
  signal ptr_deref_2004_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2004_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1898_index_0_resize_req_0 : boolean;
  signal ptr_deref_2004_load_0_ack_1 : boolean;
  signal array_obj_ref_1898_index_0_resize_ack_0 : boolean;
  signal ptr_deref_2004_load_0_req_1 : boolean;
  signal array_obj_ref_1898_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1898_index_0_rename_ack_0 : boolean;
  signal if_stmt_2063_branch_ack_0 : boolean;
  signal array_obj_ref_1898_offset_inst_req_0 : boolean;
  signal array_obj_ref_1898_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1898_base_resize_req_0 : boolean;
  signal array_obj_ref_1898_base_resize_ack_0 : boolean;
  signal binary_2087_inst_req_1 : boolean;
  signal binary_2034_inst_ack_1 : boolean;
  signal array_obj_ref_1898_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1898_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2004_load_0_ack_0 : boolean;
  signal array_obj_ref_1898_root_address_inst_req_1 : boolean;
  signal ptr_deref_2004_load_0_req_0 : boolean;
  signal array_obj_ref_1898_root_address_inst_ack_1 : boolean;
  signal binary_2034_inst_req_1 : boolean;
  signal array_obj_ref_1898_final_reg_req_0 : boolean;
  signal array_obj_ref_1898_final_reg_ack_0 : boolean;
  signal ptr_deref_1962_gather_scatter_ack_0 : boolean;
  signal binary_1944_inst_ack_1 : boolean;
  signal binary_1944_inst_req_1 : boolean;
  signal binary_1904_inst_req_0 : boolean;
  signal binary_1904_inst_ack_0 : boolean;
  signal ptr_deref_1962_gather_scatter_req_0 : boolean;
  signal binary_1904_inst_req_1 : boolean;
  signal binary_1904_inst_ack_1 : boolean;
  signal binary_1944_inst_ack_0 : boolean;
  signal ptr_deref_2004_addr_0_ack_0 : boolean;
  signal ptr_deref_1962_load_0_ack_1 : boolean;
  signal ptr_deref_2004_addr_0_req_0 : boolean;
  signal ptr_deref_1962_load_0_req_1 : boolean;
  signal binary_2044_inst_ack_1 : boolean;
  signal binary_1944_inst_req_0 : boolean;
  signal ptr_deref_2004_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2004_root_address_inst_req_0 : boolean;
  signal ptr_deref_1962_load_0_ack_0 : boolean;
  signal binary_2044_inst_req_1 : boolean;
  signal binary_2034_inst_ack_0 : boolean;
  signal array_obj_ref_1908_index_0_resize_req_0 : boolean;
  signal ptr_deref_2004_base_resize_ack_0 : boolean;
  signal array_obj_ref_1908_index_0_resize_ack_0 : boolean;
  signal ptr_deref_2004_base_resize_req_0 : boolean;
  signal array_obj_ref_1908_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1908_index_0_rename_ack_0 : boolean;
  signal if_stmt_2063_branch_ack_1 : boolean;
  signal binary_2034_inst_req_0 : boolean;
  signal array_obj_ref_1908_offset_inst_req_0 : boolean;
  signal array_obj_ref_1908_offset_inst_ack_0 : boolean;
  signal ptr_deref_1962_load_0_req_0 : boolean;
  signal array_obj_ref_1908_base_resize_req_0 : boolean;
  signal array_obj_ref_1908_base_resize_ack_0 : boolean;
  signal binary_2087_inst_ack_0 : boolean;
  signal array_obj_ref_1908_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1908_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1908_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1908_root_address_inst_ack_1 : boolean;
  signal simple_obj_ref_2070_inst_ack_0 : boolean;
  signal array_obj_ref_1908_final_reg_req_0 : boolean;
  signal binary_2000_inst_ack_1 : boolean;
  signal array_obj_ref_1908_final_reg_ack_0 : boolean;
  signal binary_2049_inst_ack_1 : boolean;
  signal binary_2049_inst_req_1 : boolean;
  signal binary_2000_inst_req_1 : boolean;
  signal binary_2000_inst_ack_0 : boolean;
  signal binary_2000_inst_req_0 : boolean;
  signal ptr_deref_1962_addr_0_ack_0 : boolean;
  signal binary_2044_inst_ack_0 : boolean;
  signal type_cast_1938_inst_ack_0 : boolean;
  signal ptr_deref_1962_addr_0_req_0 : boolean;
  signal simple_obj_ref_2070_inst_req_0 : boolean;
  signal ptr_deref_1912_base_resize_req_0 : boolean;
  signal ptr_deref_1912_base_resize_ack_0 : boolean;
  signal simple_obj_ref_2080_inst_ack_0 : boolean;
  signal type_cast_1938_inst_req_0 : boolean;
  signal ptr_deref_1912_root_address_inst_req_0 : boolean;
  signal type_cast_1994_inst_ack_0 : boolean;
  signal ptr_deref_1912_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_2080_inst_req_0 : boolean;
  signal type_cast_1994_inst_req_0 : boolean;
  signal ptr_deref_1912_addr_0_req_0 : boolean;
  signal ptr_deref_1912_addr_0_ack_0 : boolean;
  signal ptr_deref_1912_load_0_req_0 : boolean;
  signal ptr_deref_1912_load_0_ack_0 : boolean;
  signal ptr_deref_1912_load_0_req_1 : boolean;
  signal ptr_deref_1962_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1912_load_0_ack_1 : boolean;
  signal ptr_deref_1912_gather_scatter_req_0 : boolean;
  signal ptr_deref_1962_root_address_inst_req_0 : boolean;
  signal ptr_deref_1912_gather_scatter_ack_0 : boolean;
  signal binary_2055_inst_req_1 : boolean;
  signal binary_2055_inst_ack_0 : boolean;
  signal binary_2049_inst_ack_0 : boolean;
  signal ptr_deref_1990_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1990_gather_scatter_req_0 : boolean;
  signal ptr_deref_1962_base_resize_ack_0 : boolean;
  signal binary_2044_inst_req_0 : boolean;
  signal ptr_deref_1990_load_0_ack_1 : boolean;
  signal type_cast_1916_inst_req_0 : boolean;
  signal ptr_deref_1990_load_0_req_1 : boolean;
  signal type_cast_1916_inst_ack_0 : boolean;
  signal binary_2049_inst_req_0 : boolean;
  signal ptr_deref_1962_base_resize_req_0 : boolean;
  signal ptr_deref_1920_base_resize_req_0 : boolean;
  signal ptr_deref_1990_load_0_ack_0 : boolean;
  signal ptr_deref_1920_base_resize_ack_0 : boolean;
  signal ptr_deref_1934_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1990_load_0_req_0 : boolean;
  signal ptr_deref_1920_root_address_inst_req_0 : boolean;
  signal ptr_deref_1920_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1934_gather_scatter_req_0 : boolean;
  signal ptr_deref_1920_addr_0_req_0 : boolean;
  signal ptr_deref_1920_addr_0_ack_0 : boolean;
  signal ptr_deref_1934_load_0_ack_1 : boolean;
  signal ptr_deref_1920_load_0_req_0 : boolean;
  signal ptr_deref_1920_load_0_ack_0 : boolean;
  signal ptr_deref_1920_load_0_req_1 : boolean;
  signal ptr_deref_1920_load_0_ack_1 : boolean;
  signal ptr_deref_1920_gather_scatter_req_0 : boolean;
  signal ptr_deref_1920_gather_scatter_ack_0 : boolean;
  signal binary_2055_inst_req_0 : boolean;
  signal binary_2055_inst_ack_1 : boolean;
  signal ptr_deref_1934_load_0_req_1 : boolean;
  signal ptr_deref_1990_addr_0_ack_0 : boolean;
  signal ptr_deref_1990_addr_0_req_0 : boolean;
  signal binary_1958_inst_ack_1 : boolean;
  signal binary_1958_inst_req_1 : boolean;
  signal type_cast_1924_inst_req_0 : boolean;
  signal type_cast_1924_inst_ack_0 : boolean;
  signal binary_1930_inst_req_0 : boolean;
  signal binary_1930_inst_ack_0 : boolean;
  signal binary_1930_inst_req_1 : boolean;
  signal binary_1930_inst_ack_1 : boolean;
  signal simple_obj_ref_2091_inst_req_0 : boolean;
  signal simple_obj_ref_2091_inst_ack_0 : boolean;
  signal simple_obj_ref_2101_inst_req_0 : boolean;
  signal simple_obj_ref_2101_inst_ack_0 : boolean;
  signal simple_obj_ref_2110_inst_req_0 : boolean;
  signal simple_obj_ref_2110_inst_ack_0 : boolean;
  signal simple_obj_ref_2120_inst_req_0 : boolean;
  signal simple_obj_ref_2120_inst_ack_0 : boolean;
  signal phi_stmt_1816_req_1 : boolean;
  signal type_cast_1819_inst_req_0 : boolean;
  signal type_cast_1819_inst_ack_0 : boolean;
  signal phi_stmt_1816_req_0 : boolean;
  signal phi_stmt_1816_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_output_CP_7359: Block -- control-path 
    signal cp_elements: BooleanArray(518 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(489);
    cp_elements(3) <= OrReduce(cp_elements(498) & cp_elements(518));
    simple_obj_ref_2070_inst_req_0 <= cp_elements(3);
    cp_elements(4) <= simple_obj_ref_1613_inst_ack_0;
    cp_elements(5) <= cp_elements(4);
    cpelement_group_6 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(7) & cp_elements(8));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(6),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1617_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= cp_elements(5);
    cp_elements(8) <= cp_elements(5);
    cp_elements(9) <= type_cast_1617_inst_ack_0;
    cp_elements(10) <= cp_elements(5);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(10) & cp_elements(15));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1622_final_reg_req_0 <= cp_elements(11);
    cp_elements(12) <= cp_elements(9);
    array_obj_ref_1622_base_resize_req_0 <= cp_elements(12);
    cp_elements(13) <= array_obj_ref_1622_base_resize_ack_0;
    array_obj_ref_1622_root_address_inst_req_0 <= cp_elements(13);
    cp_elements(14) <= array_obj_ref_1622_root_address_inst_ack_0;
    array_obj_ref_1622_root_address_inst_req_1 <= cp_elements(14);
    cp_elements(15) <= array_obj_ref_1622_root_address_inst_ack_1;
    cp_elements(16) <= array_obj_ref_1622_final_reg_ack_0;
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(21));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1626_load_0_req_0 <= cp_elements(17);
    cp_elements(18) <= cp_elements(16);
    ptr_deref_1626_base_resize_req_0 <= cp_elements(18);
    cp_elements(19) <= ptr_deref_1626_base_resize_ack_0;
    ptr_deref_1626_root_address_inst_req_0 <= cp_elements(19);
    cp_elements(20) <= ptr_deref_1626_root_address_inst_ack_0;
    ptr_deref_1626_addr_0_req_0 <= cp_elements(20);
    cp_elements(21) <= ptr_deref_1626_addr_0_ack_0;
    cp_elements(22) <= ptr_deref_1626_load_0_ack_0;
    ptr_deref_1626_load_0_req_1 <= cp_elements(22);
    cp_elements(23) <= ptr_deref_1626_load_0_ack_1;
    ptr_deref_1626_gather_scatter_req_0 <= cp_elements(23);
    cp_elements(24) <= ptr_deref_1626_gather_scatter_ack_0;
    cpelement_group_25 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(24) & cp_elements(26));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(25),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1630_inst_req_0 <= cp_elements(25);
    cp_elements(26) <= cp_elements(5);
    cp_elements(27) <= type_cast_1630_inst_ack_0;
    cp_elements(28) <= cp_elements(5);
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(28) & cp_elements(33));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1635_final_reg_req_0 <= cp_elements(29);
    cp_elements(30) <= cp_elements(9);
    array_obj_ref_1635_base_resize_req_0 <= cp_elements(30);
    cp_elements(31) <= array_obj_ref_1635_base_resize_ack_0;
    array_obj_ref_1635_root_address_inst_req_0 <= cp_elements(31);
    cp_elements(32) <= array_obj_ref_1635_root_address_inst_ack_0;
    array_obj_ref_1635_root_address_inst_req_1 <= cp_elements(32);
    cp_elements(33) <= array_obj_ref_1635_root_address_inst_ack_1;
    cp_elements(34) <= array_obj_ref_1635_final_reg_ack_0;
    cpelement_group_35 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(34) & cp_elements(39));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(35),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1639_load_0_req_0 <= cp_elements(35);
    cp_elements(36) <= cp_elements(34);
    ptr_deref_1639_base_resize_req_0 <= cp_elements(36);
    cp_elements(37) <= ptr_deref_1639_base_resize_ack_0;
    ptr_deref_1639_root_address_inst_req_0 <= cp_elements(37);
    cp_elements(38) <= ptr_deref_1639_root_address_inst_ack_0;
    ptr_deref_1639_addr_0_req_0 <= cp_elements(38);
    cp_elements(39) <= ptr_deref_1639_addr_0_ack_0;
    cp_elements(40) <= ptr_deref_1639_load_0_ack_0;
    ptr_deref_1639_load_0_req_1 <= cp_elements(40);
    cp_elements(41) <= ptr_deref_1639_load_0_ack_1;
    ptr_deref_1639_gather_scatter_req_0 <= cp_elements(41);
    cp_elements(42) <= ptr_deref_1639_gather_scatter_ack_0;
    cpelement_group_43 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(43),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1643_inst_req_0 <= cp_elements(43);
    cp_elements(44) <= cp_elements(5);
    cp_elements(45) <= type_cast_1643_inst_ack_0;
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(47));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1649_inst_req_0 <= cp_elements(46);
    cp_elements(47) <= cp_elements(5);
    cp_elements(48) <= binary_1649_inst_ack_0;
    binary_1649_inst_req_1 <= cp_elements(48);
    cp_elements(49) <= binary_1649_inst_ack_1;
    cp_elements(50) <= cp_elements(5);
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(50) & cp_elements(55));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1654_final_reg_req_0 <= cp_elements(51);
    cp_elements(52) <= cp_elements(9);
    array_obj_ref_1654_base_resize_req_0 <= cp_elements(52);
    cp_elements(53) <= array_obj_ref_1654_base_resize_ack_0;
    array_obj_ref_1654_root_address_inst_req_0 <= cp_elements(53);
    cp_elements(54) <= array_obj_ref_1654_root_address_inst_ack_0;
    array_obj_ref_1654_root_address_inst_req_1 <= cp_elements(54);
    cp_elements(55) <= array_obj_ref_1654_root_address_inst_ack_1;
    cp_elements(56) <= array_obj_ref_1654_final_reg_ack_0;
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(61));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1658_load_0_req_0 <= cp_elements(57);
    cp_elements(58) <= cp_elements(56);
    ptr_deref_1658_base_resize_req_0 <= cp_elements(58);
    cp_elements(59) <= ptr_deref_1658_base_resize_ack_0;
    ptr_deref_1658_root_address_inst_req_0 <= cp_elements(59);
    cp_elements(60) <= ptr_deref_1658_root_address_inst_ack_0;
    ptr_deref_1658_addr_0_req_0 <= cp_elements(60);
    cp_elements(61) <= ptr_deref_1658_addr_0_ack_0;
    cp_elements(62) <= ptr_deref_1658_load_0_ack_0;
    ptr_deref_1658_load_0_req_1 <= cp_elements(62);
    cp_elements(63) <= ptr_deref_1658_load_0_ack_1;
    ptr_deref_1658_gather_scatter_req_0 <= cp_elements(63);
    cp_elements(64) <= ptr_deref_1658_gather_scatter_ack_0;
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1662_inst_req_0 <= cp_elements(65);
    cp_elements(66) <= cp_elements(5);
    cp_elements(67) <= type_cast_1662_inst_ack_0;
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(67) & cp_elements(69));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1668_inst_req_0 <= cp_elements(68);
    cp_elements(69) <= cp_elements(5);
    cp_elements(70) <= binary_1668_inst_ack_0;
    binary_1668_inst_req_1 <= cp_elements(70);
    cp_elements(71) <= binary_1668_inst_ack_1;
    cp_elements(72) <= cp_elements(5);
    cpelement_group_73 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(72) & cp_elements(77));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(73),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1673_final_reg_req_0 <= cp_elements(73);
    cp_elements(74) <= cp_elements(9);
    array_obj_ref_1673_base_resize_req_0 <= cp_elements(74);
    cp_elements(75) <= array_obj_ref_1673_base_resize_ack_0;
    array_obj_ref_1673_root_address_inst_req_0 <= cp_elements(75);
    cp_elements(76) <= array_obj_ref_1673_root_address_inst_ack_0;
    array_obj_ref_1673_root_address_inst_req_1 <= cp_elements(76);
    cp_elements(77) <= array_obj_ref_1673_root_address_inst_ack_1;
    cp_elements(78) <= array_obj_ref_1673_final_reg_ack_0;
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(83));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1677_load_0_req_0 <= cp_elements(79);
    cp_elements(80) <= cp_elements(78);
    ptr_deref_1677_base_resize_req_0 <= cp_elements(80);
    cp_elements(81) <= ptr_deref_1677_base_resize_ack_0;
    ptr_deref_1677_root_address_inst_req_0 <= cp_elements(81);
    cp_elements(82) <= ptr_deref_1677_root_address_inst_ack_0;
    ptr_deref_1677_addr_0_req_0 <= cp_elements(82);
    cp_elements(83) <= ptr_deref_1677_addr_0_ack_0;
    cp_elements(84) <= ptr_deref_1677_load_0_ack_0;
    ptr_deref_1677_load_0_req_1 <= cp_elements(84);
    cp_elements(85) <= ptr_deref_1677_load_0_ack_1;
    ptr_deref_1677_gather_scatter_req_0 <= cp_elements(85);
    cp_elements(86) <= ptr_deref_1677_gather_scatter_ack_0;
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(86) & cp_elements(88));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1681_inst_req_0 <= cp_elements(87);
    cp_elements(88) <= cp_elements(5);
    cp_elements(89) <= type_cast_1681_inst_ack_0;
    cpelement_group_90 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(91));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(90),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1687_inst_req_0 <= cp_elements(90);
    cp_elements(91) <= cp_elements(5);
    cp_elements(92) <= binary_1687_inst_ack_0;
    binary_1687_inst_req_1 <= cp_elements(92);
    cp_elements(93) <= binary_1687_inst_ack_1;
    cp_elements(94) <= cp_elements(5);
    cpelement_group_95 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(94) & cp_elements(99));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(95),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1692_final_reg_req_0 <= cp_elements(95);
    cp_elements(96) <= cp_elements(9);
    array_obj_ref_1692_base_resize_req_0 <= cp_elements(96);
    cp_elements(97) <= array_obj_ref_1692_base_resize_ack_0;
    array_obj_ref_1692_root_address_inst_req_0 <= cp_elements(97);
    cp_elements(98) <= array_obj_ref_1692_root_address_inst_ack_0;
    array_obj_ref_1692_root_address_inst_req_1 <= cp_elements(98);
    cp_elements(99) <= array_obj_ref_1692_root_address_inst_ack_1;
    cp_elements(100) <= array_obj_ref_1692_final_reg_ack_0;
    cpelement_group_101 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(100) & cp_elements(105));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(101),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1696_load_0_req_0 <= cp_elements(101);
    cp_elements(102) <= cp_elements(100);
    ptr_deref_1696_base_resize_req_0 <= cp_elements(102);
    cp_elements(103) <= ptr_deref_1696_base_resize_ack_0;
    ptr_deref_1696_root_address_inst_req_0 <= cp_elements(103);
    cp_elements(104) <= ptr_deref_1696_root_address_inst_ack_0;
    ptr_deref_1696_addr_0_req_0 <= cp_elements(104);
    cp_elements(105) <= ptr_deref_1696_addr_0_ack_0;
    cp_elements(106) <= ptr_deref_1696_load_0_ack_0;
    ptr_deref_1696_load_0_req_1 <= cp_elements(106);
    cp_elements(107) <= ptr_deref_1696_load_0_ack_1;
    ptr_deref_1696_gather_scatter_req_0 <= cp_elements(107);
    cp_elements(108) <= ptr_deref_1696_gather_scatter_ack_0;
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(108) & cp_elements(110));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1700_inst_req_0 <= cp_elements(109);
    cp_elements(110) <= cp_elements(5);
    cp_elements(111) <= type_cast_1700_inst_ack_0;
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(111) & cp_elements(113));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1706_inst_req_0 <= cp_elements(112);
    cp_elements(113) <= cp_elements(5);
    cp_elements(114) <= binary_1706_inst_ack_0;
    binary_1706_inst_req_1 <= cp_elements(114);
    cp_elements(115) <= binary_1706_inst_ack_1;
    cp_elements(116) <= cp_elements(5);
    cpelement_group_117 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(116) & cp_elements(121));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(117),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1711_final_reg_req_0 <= cp_elements(117);
    cp_elements(118) <= cp_elements(9);
    array_obj_ref_1711_base_resize_req_0 <= cp_elements(118);
    cp_elements(119) <= array_obj_ref_1711_base_resize_ack_0;
    array_obj_ref_1711_root_address_inst_req_0 <= cp_elements(119);
    cp_elements(120) <= array_obj_ref_1711_root_address_inst_ack_0;
    array_obj_ref_1711_root_address_inst_req_1 <= cp_elements(120);
    cp_elements(121) <= array_obj_ref_1711_root_address_inst_ack_1;
    cp_elements(122) <= array_obj_ref_1711_final_reg_ack_0;
    cpelement_group_123 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(122) & cp_elements(127));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(123),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1715_load_0_req_0 <= cp_elements(123);
    cp_elements(124) <= cp_elements(122);
    ptr_deref_1715_base_resize_req_0 <= cp_elements(124);
    cp_elements(125) <= ptr_deref_1715_base_resize_ack_0;
    ptr_deref_1715_root_address_inst_req_0 <= cp_elements(125);
    cp_elements(126) <= ptr_deref_1715_root_address_inst_ack_0;
    ptr_deref_1715_addr_0_req_0 <= cp_elements(126);
    cp_elements(127) <= ptr_deref_1715_addr_0_ack_0;
    cp_elements(128) <= ptr_deref_1715_load_0_ack_0;
    ptr_deref_1715_load_0_req_1 <= cp_elements(128);
    cp_elements(129) <= ptr_deref_1715_load_0_ack_1;
    ptr_deref_1715_gather_scatter_req_0 <= cp_elements(129);
    cp_elements(130) <= ptr_deref_1715_gather_scatter_ack_0;
    cpelement_group_131 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(130) & cp_elements(132));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(131),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1719_inst_req_0 <= cp_elements(131);
    cp_elements(132) <= cp_elements(5);
    cp_elements(133) <= type_cast_1719_inst_ack_0;
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(133) & cp_elements(135));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1725_inst_req_0 <= cp_elements(134);
    cp_elements(135) <= cp_elements(5);
    cp_elements(136) <= binary_1725_inst_ack_0;
    binary_1725_inst_req_1 <= cp_elements(136);
    cp_elements(137) <= binary_1725_inst_ack_1;
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(143));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1729_load_0_req_0 <= cp_elements(138);
    cp_elements(139) <= cp_elements(9);
    cp_elements(140) <= cp_elements(139);
    ptr_deref_1729_base_resize_req_0 <= cp_elements(140);
    cp_elements(141) <= ptr_deref_1729_base_resize_ack_0;
    ptr_deref_1729_root_address_inst_req_0 <= cp_elements(141);
    cp_elements(142) <= ptr_deref_1729_root_address_inst_ack_0;
    ptr_deref_1729_addr_0_req_0 <= cp_elements(142);
    cp_elements(143) <= ptr_deref_1729_addr_0_ack_0;
    cp_elements(144) <= ptr_deref_1729_load_0_ack_0;
    ptr_deref_1729_load_0_req_1 <= cp_elements(144);
    cp_elements(145) <= ptr_deref_1729_load_0_ack_1;
    ptr_deref_1729_gather_scatter_req_0 <= cp_elements(145);
    cp_elements(146) <= ptr_deref_1729_gather_scatter_ack_0;
    cpelement_group_147 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(146) & cp_elements(148));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1733_inst_req_0 <= cp_elements(147);
    cp_elements(148) <= cp_elements(5);
    cp_elements(149) <= type_cast_1733_inst_ack_0;
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(151));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1739_inst_req_0 <= cp_elements(150);
    cp_elements(151) <= cp_elements(5);
    cp_elements(152) <= binary_1739_inst_ack_0;
    binary_1739_inst_req_1 <= cp_elements(152);
    cp_elements(153) <= binary_1739_inst_ack_1;
    cp_elements(154) <= cp_elements(5);
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(154) & cp_elements(159));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1744_final_reg_req_0 <= cp_elements(155);
    cp_elements(156) <= cp_elements(9);
    array_obj_ref_1744_base_resize_req_0 <= cp_elements(156);
    cp_elements(157) <= array_obj_ref_1744_base_resize_ack_0;
    array_obj_ref_1744_root_address_inst_req_0 <= cp_elements(157);
    cp_elements(158) <= array_obj_ref_1744_root_address_inst_ack_0;
    array_obj_ref_1744_root_address_inst_req_1 <= cp_elements(158);
    cp_elements(159) <= array_obj_ref_1744_root_address_inst_ack_1;
    cp_elements(160) <= array_obj_ref_1744_final_reg_ack_0;
    cpelement_group_161 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(160) & cp_elements(165));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(161),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1748_load_0_req_0 <= cp_elements(161);
    cp_elements(162) <= cp_elements(160);
    ptr_deref_1748_base_resize_req_0 <= cp_elements(162);
    cp_elements(163) <= ptr_deref_1748_base_resize_ack_0;
    ptr_deref_1748_root_address_inst_req_0 <= cp_elements(163);
    cp_elements(164) <= ptr_deref_1748_root_address_inst_ack_0;
    ptr_deref_1748_addr_0_req_0 <= cp_elements(164);
    cp_elements(165) <= ptr_deref_1748_addr_0_ack_0;
    cp_elements(166) <= ptr_deref_1748_load_0_ack_0;
    ptr_deref_1748_load_0_req_1 <= cp_elements(166);
    cp_elements(167) <= ptr_deref_1748_load_0_ack_1;
    ptr_deref_1748_gather_scatter_req_0 <= cp_elements(167);
    cp_elements(168) <= ptr_deref_1748_gather_scatter_ack_0;
    cpelement_group_169 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(168) & cp_elements(170));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(169),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1752_inst_req_0 <= cp_elements(169);
    cp_elements(170) <= cp_elements(5);
    cp_elements(171) <= type_cast_1752_inst_ack_0;
    cpelement_group_172 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(171) & cp_elements(173));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(172),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1758_inst_req_0 <= cp_elements(172);
    cp_elements(173) <= cp_elements(5);
    cp_elements(174) <= binary_1758_inst_ack_0;
    binary_1758_inst_req_1 <= cp_elements(174);
    cp_elements(175) <= binary_1758_inst_ack_1;
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(49) & cp_elements(177));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1763_inst_req_0 <= cp_elements(176);
    cp_elements(177) <= cp_elements(5);
    cp_elements(178) <= binary_1763_inst_ack_0;
    binary_1763_inst_req_1 <= cp_elements(178);
    cp_elements(179) <= binary_1763_inst_ack_1;
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(179) & cp_elements(181));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1768_inst_req_0 <= cp_elements(180);
    cp_elements(181) <= cp_elements(5);
    cp_elements(182) <= binary_1768_inst_ack_0;
    binary_1768_inst_req_1 <= cp_elements(182);
    cp_elements(183) <= binary_1768_inst_ack_1;
    cpelement_group_184 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(183) & cp_elements(185));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(184),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1773_inst_req_0 <= cp_elements(184);
    cp_elements(185) <= cp_elements(5);
    cp_elements(186) <= binary_1773_inst_ack_0;
    binary_1773_inst_req_1 <= cp_elements(186);
    cp_elements(187) <= binary_1773_inst_ack_1;
    cpelement_group_188 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(115) & cp_elements(187) & cp_elements(189));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(188),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1778_inst_req_0 <= cp_elements(188);
    cp_elements(189) <= cp_elements(5);
    cp_elements(190) <= binary_1778_inst_ack_0;
    binary_1778_inst_req_1 <= cp_elements(190);
    cp_elements(191) <= binary_1778_inst_ack_1;
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1783_inst_req_0 <= cp_elements(192);
    cp_elements(193) <= cp_elements(5);
    cp_elements(194) <= binary_1783_inst_ack_0;
    binary_1783_inst_req_1 <= cp_elements(194);
    cp_elements(195) <= binary_1783_inst_ack_1;
    cpelement_group_196 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(153) & cp_elements(195) & cp_elements(197));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(196),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1788_inst_req_0 <= cp_elements(196);
    cp_elements(197) <= cp_elements(5);
    cp_elements(198) <= binary_1788_inst_ack_0;
    binary_1788_inst_req_1 <= cp_elements(198);
    cp_elements(199) <= binary_1788_inst_ack_1;
    cpelement_group_200 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(199) & cp_elements(201));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(200),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1793_inst_req_0 <= cp_elements(200);
    cp_elements(201) <= cp_elements(5);
    cp_elements(202) <= binary_1793_inst_ack_0;
    binary_1793_inst_req_1 <= cp_elements(202);
    cp_elements(203) <= binary_1793_inst_ack_1;
    simple_obj_ref_1801_inst_req_0 <= cp_elements(203);
    cp_elements(204) <= simple_obj_ref_1801_inst_ack_0;
    simple_obj_ref_1811_inst_req_0 <= cp_elements(204);
    cp_elements(205) <= simple_obj_ref_1811_inst_ack_0;
    phi_stmt_1816_req_1 <= cp_elements(205);
    cp_elements(206) <= cp_elements(516);
    cpelement_group_207 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(208) & cp_elements(209));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(207),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1828_inst_req_0 <= cp_elements(207);
    cp_elements(208) <= cp_elements(206);
    cp_elements(209) <= cp_elements(206);
    cp_elements(210) <= binary_1828_inst_ack_0;
    binary_1828_inst_req_1 <= cp_elements(210);
    cp_elements(211) <= binary_1828_inst_ack_1;
    cpelement_group_212 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(213) & cp_elements(214));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(212),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1834_inst_req_0 <= cp_elements(212);
    cp_elements(213) <= cp_elements(206);
    cp_elements(214) <= cp_elements(211);
    cp_elements(215) <= binary_1834_inst_ack_0;
    binary_1834_inst_req_1 <= cp_elements(215);
    cp_elements(216) <= binary_1834_inst_ack_1;
    array_obj_ref_1838_index_0_resize_req_0 <= cp_elements(216);
    cp_elements(217) <= cp_elements(206);
    cpelement_group_218 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(217) & cp_elements(226));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(218),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1838_final_reg_req_0 <= cp_elements(218);
    cp_elements(219) <= cp_elements(206);
    array_obj_ref_1838_base_resize_req_0 <= cp_elements(219);
    cp_elements(220) <= array_obj_ref_1838_index_0_resize_ack_0;
    array_obj_ref_1838_index_0_rename_req_0 <= cp_elements(220);
    cp_elements(221) <= array_obj_ref_1838_index_0_rename_ack_0;
    array_obj_ref_1838_offset_inst_req_0 <= cp_elements(221);
    cp_elements(222) <= array_obj_ref_1838_offset_inst_ack_0;
    cp_elements(223) <= array_obj_ref_1838_base_resize_ack_0;
    cpelement_group_224 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(222) & cp_elements(223));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(224),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1838_root_address_inst_req_0 <= cp_elements(224);
    cp_elements(225) <= array_obj_ref_1838_root_address_inst_ack_0;
    array_obj_ref_1838_root_address_inst_req_1 <= cp_elements(225);
    cp_elements(226) <= array_obj_ref_1838_root_address_inst_ack_1;
    cp_elements(227) <= array_obj_ref_1838_final_reg_ack_0;
    cpelement_group_228 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(229) & cp_elements(230));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(228),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1844_inst_req_0 <= cp_elements(228);
    cp_elements(229) <= cp_elements(206);
    cp_elements(230) <= cp_elements(211);
    cp_elements(231) <= binary_1844_inst_ack_0;
    binary_1844_inst_req_1 <= cp_elements(231);
    cp_elements(232) <= binary_1844_inst_ack_1;
    array_obj_ref_1848_index_0_resize_req_0 <= cp_elements(232);
    cp_elements(233) <= cp_elements(206);
    cpelement_group_234 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(233) & cp_elements(242));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(234),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1848_final_reg_req_0 <= cp_elements(234);
    cp_elements(235) <= cp_elements(206);
    array_obj_ref_1848_base_resize_req_0 <= cp_elements(235);
    cp_elements(236) <= array_obj_ref_1848_index_0_resize_ack_0;
    array_obj_ref_1848_index_0_rename_req_0 <= cp_elements(236);
    cp_elements(237) <= array_obj_ref_1848_index_0_rename_ack_0;
    array_obj_ref_1848_offset_inst_req_0 <= cp_elements(237);
    cp_elements(238) <= array_obj_ref_1848_offset_inst_ack_0;
    cp_elements(239) <= array_obj_ref_1848_base_resize_ack_0;
    cpelement_group_240 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(239));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(240),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1848_root_address_inst_req_0 <= cp_elements(240);
    cp_elements(241) <= array_obj_ref_1848_root_address_inst_ack_0;
    array_obj_ref_1848_root_address_inst_req_1 <= cp_elements(241);
    cp_elements(242) <= array_obj_ref_1848_root_address_inst_ack_1;
    cp_elements(243) <= array_obj_ref_1848_final_reg_ack_0;
    cpelement_group_244 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(246));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(244),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1854_inst_req_0 <= cp_elements(244);
    cp_elements(245) <= cp_elements(206);
    cp_elements(246) <= cp_elements(211);
    cp_elements(247) <= binary_1854_inst_ack_0;
    binary_1854_inst_req_1 <= cp_elements(247);
    cp_elements(248) <= binary_1854_inst_ack_1;
    array_obj_ref_1858_index_0_resize_req_0 <= cp_elements(248);
    cp_elements(249) <= cp_elements(206);
    cpelement_group_250 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(249) & cp_elements(258));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(250),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1858_final_reg_req_0 <= cp_elements(250);
    cp_elements(251) <= cp_elements(206);
    array_obj_ref_1858_base_resize_req_0 <= cp_elements(251);
    cp_elements(252) <= array_obj_ref_1858_index_0_resize_ack_0;
    array_obj_ref_1858_index_0_rename_req_0 <= cp_elements(252);
    cp_elements(253) <= array_obj_ref_1858_index_0_rename_ack_0;
    array_obj_ref_1858_offset_inst_req_0 <= cp_elements(253);
    cp_elements(254) <= array_obj_ref_1858_offset_inst_ack_0;
    cp_elements(255) <= array_obj_ref_1858_base_resize_ack_0;
    cpelement_group_256 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(255));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(256),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1858_root_address_inst_req_0 <= cp_elements(256);
    cp_elements(257) <= array_obj_ref_1858_root_address_inst_ack_0;
    array_obj_ref_1858_root_address_inst_req_1 <= cp_elements(257);
    cp_elements(258) <= array_obj_ref_1858_root_address_inst_ack_1;
    cp_elements(259) <= array_obj_ref_1858_final_reg_ack_0;
    cpelement_group_260 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(261) & cp_elements(262));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(260),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1864_inst_req_0 <= cp_elements(260);
    cp_elements(261) <= cp_elements(206);
    cp_elements(262) <= cp_elements(211);
    cp_elements(263) <= binary_1864_inst_ack_0;
    binary_1864_inst_req_1 <= cp_elements(263);
    cp_elements(264) <= binary_1864_inst_ack_1;
    array_obj_ref_1868_index_0_resize_req_0 <= cp_elements(264);
    cp_elements(265) <= cp_elements(206);
    cpelement_group_266 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(265) & cp_elements(274));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(266),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1868_final_reg_req_0 <= cp_elements(266);
    cp_elements(267) <= cp_elements(206);
    array_obj_ref_1868_base_resize_req_0 <= cp_elements(267);
    cp_elements(268) <= array_obj_ref_1868_index_0_resize_ack_0;
    array_obj_ref_1868_index_0_rename_req_0 <= cp_elements(268);
    cp_elements(269) <= array_obj_ref_1868_index_0_rename_ack_0;
    array_obj_ref_1868_offset_inst_req_0 <= cp_elements(269);
    cp_elements(270) <= array_obj_ref_1868_offset_inst_ack_0;
    cp_elements(271) <= array_obj_ref_1868_base_resize_ack_0;
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(270) & cp_elements(271));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1868_root_address_inst_req_0 <= cp_elements(272);
    cp_elements(273) <= array_obj_ref_1868_root_address_inst_ack_0;
    array_obj_ref_1868_root_address_inst_req_1 <= cp_elements(273);
    cp_elements(274) <= array_obj_ref_1868_root_address_inst_ack_1;
    cp_elements(275) <= array_obj_ref_1868_final_reg_ack_0;
    cpelement_group_276 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(277) & cp_elements(278));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(276),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1874_inst_req_0 <= cp_elements(276);
    cp_elements(277) <= cp_elements(206);
    cp_elements(278) <= cp_elements(211);
    cp_elements(279) <= binary_1874_inst_ack_0;
    binary_1874_inst_req_1 <= cp_elements(279);
    cp_elements(280) <= binary_1874_inst_ack_1;
    array_obj_ref_1878_index_0_resize_req_0 <= cp_elements(280);
    cp_elements(281) <= cp_elements(206);
    cpelement_group_282 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(281) & cp_elements(290));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(282),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1878_final_reg_req_0 <= cp_elements(282);
    cp_elements(283) <= cp_elements(206);
    array_obj_ref_1878_base_resize_req_0 <= cp_elements(283);
    cp_elements(284) <= array_obj_ref_1878_index_0_resize_ack_0;
    array_obj_ref_1878_index_0_rename_req_0 <= cp_elements(284);
    cp_elements(285) <= array_obj_ref_1878_index_0_rename_ack_0;
    array_obj_ref_1878_offset_inst_req_0 <= cp_elements(285);
    cp_elements(286) <= array_obj_ref_1878_offset_inst_ack_0;
    cp_elements(287) <= array_obj_ref_1878_base_resize_ack_0;
    cpelement_group_288 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(286) & cp_elements(287));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(288),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1878_root_address_inst_req_0 <= cp_elements(288);
    cp_elements(289) <= array_obj_ref_1878_root_address_inst_ack_0;
    array_obj_ref_1878_root_address_inst_req_1 <= cp_elements(289);
    cp_elements(290) <= array_obj_ref_1878_root_address_inst_ack_1;
    cp_elements(291) <= array_obj_ref_1878_final_reg_ack_0;
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(293) & cp_elements(294));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1884_inst_req_0 <= cp_elements(292);
    cp_elements(293) <= cp_elements(206);
    cp_elements(294) <= cp_elements(211);
    cp_elements(295) <= binary_1884_inst_ack_0;
    binary_1884_inst_req_1 <= cp_elements(295);
    cp_elements(296) <= binary_1884_inst_ack_1;
    array_obj_ref_1888_index_0_resize_req_0 <= cp_elements(296);
    cp_elements(297) <= cp_elements(206);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(297) & cp_elements(306));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1888_final_reg_req_0 <= cp_elements(298);
    cp_elements(299) <= cp_elements(206);
    array_obj_ref_1888_base_resize_req_0 <= cp_elements(299);
    cp_elements(300) <= array_obj_ref_1888_index_0_resize_ack_0;
    array_obj_ref_1888_index_0_rename_req_0 <= cp_elements(300);
    cp_elements(301) <= array_obj_ref_1888_index_0_rename_ack_0;
    array_obj_ref_1888_offset_inst_req_0 <= cp_elements(301);
    cp_elements(302) <= array_obj_ref_1888_offset_inst_ack_0;
    cp_elements(303) <= array_obj_ref_1888_base_resize_ack_0;
    cpelement_group_304 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(302) & cp_elements(303));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(304),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1888_root_address_inst_req_0 <= cp_elements(304);
    cp_elements(305) <= array_obj_ref_1888_root_address_inst_ack_0;
    array_obj_ref_1888_root_address_inst_req_1 <= cp_elements(305);
    cp_elements(306) <= array_obj_ref_1888_root_address_inst_ack_1;
    cp_elements(307) <= array_obj_ref_1888_final_reg_ack_0;
    cpelement_group_308 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(309) & cp_elements(310));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1894_inst_req_0 <= cp_elements(308);
    cp_elements(309) <= cp_elements(206);
    cp_elements(310) <= cp_elements(211);
    cp_elements(311) <= binary_1894_inst_ack_0;
    binary_1894_inst_req_1 <= cp_elements(311);
    cp_elements(312) <= binary_1894_inst_ack_1;
    array_obj_ref_1898_index_0_resize_req_0 <= cp_elements(312);
    cp_elements(313) <= cp_elements(206);
    cpelement_group_314 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(313) & cp_elements(322));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(314),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1898_final_reg_req_0 <= cp_elements(314);
    cp_elements(315) <= cp_elements(206);
    array_obj_ref_1898_base_resize_req_0 <= cp_elements(315);
    cp_elements(316) <= array_obj_ref_1898_index_0_resize_ack_0;
    array_obj_ref_1898_index_0_rename_req_0 <= cp_elements(316);
    cp_elements(317) <= array_obj_ref_1898_index_0_rename_ack_0;
    array_obj_ref_1898_offset_inst_req_0 <= cp_elements(317);
    cp_elements(318) <= array_obj_ref_1898_offset_inst_ack_0;
    cp_elements(319) <= array_obj_ref_1898_base_resize_ack_0;
    cpelement_group_320 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(318) & cp_elements(319));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(320),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1898_root_address_inst_req_0 <= cp_elements(320);
    cp_elements(321) <= array_obj_ref_1898_root_address_inst_ack_0;
    array_obj_ref_1898_root_address_inst_req_1 <= cp_elements(321);
    cp_elements(322) <= array_obj_ref_1898_root_address_inst_ack_1;
    cp_elements(323) <= array_obj_ref_1898_final_reg_ack_0;
    cpelement_group_324 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(325) & cp_elements(326));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(324),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1904_inst_req_0 <= cp_elements(324);
    cp_elements(325) <= cp_elements(206);
    cp_elements(326) <= cp_elements(211);
    cp_elements(327) <= binary_1904_inst_ack_0;
    binary_1904_inst_req_1 <= cp_elements(327);
    cp_elements(328) <= binary_1904_inst_ack_1;
    array_obj_ref_1908_index_0_resize_req_0 <= cp_elements(328);
    cp_elements(329) <= cp_elements(206);
    cpelement_group_330 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(329) & cp_elements(338));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(330),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1908_final_reg_req_0 <= cp_elements(330);
    cp_elements(331) <= cp_elements(206);
    array_obj_ref_1908_base_resize_req_0 <= cp_elements(331);
    cp_elements(332) <= array_obj_ref_1908_index_0_resize_ack_0;
    array_obj_ref_1908_index_0_rename_req_0 <= cp_elements(332);
    cp_elements(333) <= array_obj_ref_1908_index_0_rename_ack_0;
    array_obj_ref_1908_offset_inst_req_0 <= cp_elements(333);
    cp_elements(334) <= array_obj_ref_1908_offset_inst_ack_0;
    cp_elements(335) <= array_obj_ref_1908_base_resize_ack_0;
    cpelement_group_336 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(334) & cp_elements(335));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(336),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1908_root_address_inst_req_0 <= cp_elements(336);
    cp_elements(337) <= array_obj_ref_1908_root_address_inst_ack_0;
    array_obj_ref_1908_root_address_inst_req_1 <= cp_elements(337);
    cp_elements(338) <= array_obj_ref_1908_root_address_inst_ack_1;
    cp_elements(339) <= array_obj_ref_1908_final_reg_ack_0;
    cpelement_group_340 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(339) & cp_elements(344));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(340),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1912_load_0_req_0 <= cp_elements(340);
    cp_elements(341) <= cp_elements(339);
    ptr_deref_1912_base_resize_req_0 <= cp_elements(341);
    cp_elements(342) <= ptr_deref_1912_base_resize_ack_0;
    ptr_deref_1912_root_address_inst_req_0 <= cp_elements(342);
    cp_elements(343) <= ptr_deref_1912_root_address_inst_ack_0;
    ptr_deref_1912_addr_0_req_0 <= cp_elements(343);
    cp_elements(344) <= ptr_deref_1912_addr_0_ack_0;
    cp_elements(345) <= ptr_deref_1912_load_0_ack_0;
    ptr_deref_1912_load_0_req_1 <= cp_elements(345);
    cp_elements(346) <= ptr_deref_1912_load_0_ack_1;
    ptr_deref_1912_gather_scatter_req_0 <= cp_elements(346);
    cp_elements(347) <= ptr_deref_1912_gather_scatter_ack_0;
    cpelement_group_348 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(347) & cp_elements(349));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(348),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1916_inst_req_0 <= cp_elements(348);
    cp_elements(349) <= cp_elements(206);
    cp_elements(350) <= type_cast_1916_inst_ack_0;
    cpelement_group_351 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(323) & cp_elements(355));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(351),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1920_load_0_req_0 <= cp_elements(351);
    cp_elements(352) <= cp_elements(323);
    ptr_deref_1920_base_resize_req_0 <= cp_elements(352);
    cp_elements(353) <= ptr_deref_1920_base_resize_ack_0;
    ptr_deref_1920_root_address_inst_req_0 <= cp_elements(353);
    cp_elements(354) <= ptr_deref_1920_root_address_inst_ack_0;
    ptr_deref_1920_addr_0_req_0 <= cp_elements(354);
    cp_elements(355) <= ptr_deref_1920_addr_0_ack_0;
    cp_elements(356) <= ptr_deref_1920_load_0_ack_0;
    ptr_deref_1920_load_0_req_1 <= cp_elements(356);
    cp_elements(357) <= ptr_deref_1920_load_0_ack_1;
    ptr_deref_1920_gather_scatter_req_0 <= cp_elements(357);
    cp_elements(358) <= ptr_deref_1920_gather_scatter_ack_0;
    cpelement_group_359 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(358) & cp_elements(360));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(359),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1924_inst_req_0 <= cp_elements(359);
    cp_elements(360) <= cp_elements(206);
    cp_elements(361) <= type_cast_1924_inst_ack_0;
    cpelement_group_362 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(361) & cp_elements(363));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(362),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1930_inst_req_0 <= cp_elements(362);
    cp_elements(363) <= cp_elements(206);
    cp_elements(364) <= binary_1930_inst_ack_0;
    binary_1930_inst_req_1 <= cp_elements(364);
    cp_elements(365) <= binary_1930_inst_ack_1;
    cpelement_group_366 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(307) & cp_elements(370));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(366),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1934_load_0_req_0 <= cp_elements(366);
    cp_elements(367) <= cp_elements(307);
    ptr_deref_1934_base_resize_req_0 <= cp_elements(367);
    cp_elements(368) <= ptr_deref_1934_base_resize_ack_0;
    ptr_deref_1934_root_address_inst_req_0 <= cp_elements(368);
    cp_elements(369) <= ptr_deref_1934_root_address_inst_ack_0;
    ptr_deref_1934_addr_0_req_0 <= cp_elements(369);
    cp_elements(370) <= ptr_deref_1934_addr_0_ack_0;
    cp_elements(371) <= ptr_deref_1934_load_0_ack_0;
    ptr_deref_1934_load_0_req_1 <= cp_elements(371);
    cp_elements(372) <= ptr_deref_1934_load_0_ack_1;
    ptr_deref_1934_gather_scatter_req_0 <= cp_elements(372);
    cp_elements(373) <= ptr_deref_1934_gather_scatter_ack_0;
    cpelement_group_374 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(373) & cp_elements(375));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(374),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1938_inst_req_0 <= cp_elements(374);
    cp_elements(375) <= cp_elements(206);
    cp_elements(376) <= type_cast_1938_inst_ack_0;
    cpelement_group_377 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(376) & cp_elements(378));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(377),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1944_inst_req_0 <= cp_elements(377);
    cp_elements(378) <= cp_elements(206);
    cp_elements(379) <= binary_1944_inst_ack_0;
    binary_1944_inst_req_1 <= cp_elements(379);
    cp_elements(380) <= binary_1944_inst_ack_1;
    cpelement_group_381 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(385));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(381),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1948_load_0_req_0 <= cp_elements(381);
    cp_elements(382) <= cp_elements(291);
    ptr_deref_1948_base_resize_req_0 <= cp_elements(382);
    cp_elements(383) <= ptr_deref_1948_base_resize_ack_0;
    ptr_deref_1948_root_address_inst_req_0 <= cp_elements(383);
    cp_elements(384) <= ptr_deref_1948_root_address_inst_ack_0;
    ptr_deref_1948_addr_0_req_0 <= cp_elements(384);
    cp_elements(385) <= ptr_deref_1948_addr_0_ack_0;
    cp_elements(386) <= ptr_deref_1948_load_0_ack_0;
    ptr_deref_1948_load_0_req_1 <= cp_elements(386);
    cp_elements(387) <= ptr_deref_1948_load_0_ack_1;
    ptr_deref_1948_gather_scatter_req_0 <= cp_elements(387);
    cp_elements(388) <= ptr_deref_1948_gather_scatter_ack_0;
    cpelement_group_389 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(388) & cp_elements(390));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(389),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1952_inst_req_0 <= cp_elements(389);
    cp_elements(390) <= cp_elements(206);
    cp_elements(391) <= type_cast_1952_inst_ack_0;
    cpelement_group_392 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(391) & cp_elements(393));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(392),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1958_inst_req_0 <= cp_elements(392);
    cp_elements(393) <= cp_elements(206);
    cp_elements(394) <= binary_1958_inst_ack_0;
    binary_1958_inst_req_1 <= cp_elements(394);
    cp_elements(395) <= binary_1958_inst_ack_1;
    cpelement_group_396 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(275) & cp_elements(400));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(396),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1962_load_0_req_0 <= cp_elements(396);
    cp_elements(397) <= cp_elements(275);
    ptr_deref_1962_base_resize_req_0 <= cp_elements(397);
    cp_elements(398) <= ptr_deref_1962_base_resize_ack_0;
    ptr_deref_1962_root_address_inst_req_0 <= cp_elements(398);
    cp_elements(399) <= ptr_deref_1962_root_address_inst_ack_0;
    ptr_deref_1962_addr_0_req_0 <= cp_elements(399);
    cp_elements(400) <= ptr_deref_1962_addr_0_ack_0;
    cp_elements(401) <= ptr_deref_1962_load_0_ack_0;
    ptr_deref_1962_load_0_req_1 <= cp_elements(401);
    cp_elements(402) <= ptr_deref_1962_load_0_ack_1;
    ptr_deref_1962_gather_scatter_req_0 <= cp_elements(402);
    cp_elements(403) <= ptr_deref_1962_gather_scatter_ack_0;
    cpelement_group_404 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(403) & cp_elements(405));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(404),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1966_inst_req_0 <= cp_elements(404);
    cp_elements(405) <= cp_elements(206);
    cp_elements(406) <= type_cast_1966_inst_ack_0;
    cpelement_group_407 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(406) & cp_elements(408));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(407),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1972_inst_req_0 <= cp_elements(407);
    cp_elements(408) <= cp_elements(206);
    cp_elements(409) <= binary_1972_inst_ack_0;
    binary_1972_inst_req_1 <= cp_elements(409);
    cp_elements(410) <= binary_1972_inst_ack_1;
    cpelement_group_411 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(259) & cp_elements(415));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(411),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1976_load_0_req_0 <= cp_elements(411);
    cp_elements(412) <= cp_elements(259);
    ptr_deref_1976_base_resize_req_0 <= cp_elements(412);
    cp_elements(413) <= ptr_deref_1976_base_resize_ack_0;
    ptr_deref_1976_root_address_inst_req_0 <= cp_elements(413);
    cp_elements(414) <= ptr_deref_1976_root_address_inst_ack_0;
    ptr_deref_1976_addr_0_req_0 <= cp_elements(414);
    cp_elements(415) <= ptr_deref_1976_addr_0_ack_0;
    cp_elements(416) <= ptr_deref_1976_load_0_ack_0;
    ptr_deref_1976_load_0_req_1 <= cp_elements(416);
    cp_elements(417) <= ptr_deref_1976_load_0_ack_1;
    ptr_deref_1976_gather_scatter_req_0 <= cp_elements(417);
    cp_elements(418) <= ptr_deref_1976_gather_scatter_ack_0;
    cpelement_group_419 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(418) & cp_elements(420));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(419),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1980_inst_req_0 <= cp_elements(419);
    cp_elements(420) <= cp_elements(206);
    cp_elements(421) <= type_cast_1980_inst_ack_0;
    cpelement_group_422 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(421) & cp_elements(423));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(422),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1986_inst_req_0 <= cp_elements(422);
    cp_elements(423) <= cp_elements(206);
    cp_elements(424) <= binary_1986_inst_ack_0;
    binary_1986_inst_req_1 <= cp_elements(424);
    cp_elements(425) <= binary_1986_inst_ack_1;
    cpelement_group_426 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(243) & cp_elements(430));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(426),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1990_load_0_req_0 <= cp_elements(426);
    cp_elements(427) <= cp_elements(243);
    ptr_deref_1990_base_resize_req_0 <= cp_elements(427);
    cp_elements(428) <= ptr_deref_1990_base_resize_ack_0;
    ptr_deref_1990_root_address_inst_req_0 <= cp_elements(428);
    cp_elements(429) <= ptr_deref_1990_root_address_inst_ack_0;
    ptr_deref_1990_addr_0_req_0 <= cp_elements(429);
    cp_elements(430) <= ptr_deref_1990_addr_0_ack_0;
    cp_elements(431) <= ptr_deref_1990_load_0_ack_0;
    ptr_deref_1990_load_0_req_1 <= cp_elements(431);
    cp_elements(432) <= ptr_deref_1990_load_0_ack_1;
    ptr_deref_1990_gather_scatter_req_0 <= cp_elements(432);
    cp_elements(433) <= ptr_deref_1990_gather_scatter_ack_0;
    cpelement_group_434 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(433) & cp_elements(435));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(434),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1994_inst_req_0 <= cp_elements(434);
    cp_elements(435) <= cp_elements(206);
    cp_elements(436) <= type_cast_1994_inst_ack_0;
    cpelement_group_437 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(436) & cp_elements(438));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(437),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2000_inst_req_0 <= cp_elements(437);
    cp_elements(438) <= cp_elements(206);
    cp_elements(439) <= binary_2000_inst_ack_0;
    binary_2000_inst_req_1 <= cp_elements(439);
    cp_elements(440) <= binary_2000_inst_ack_1;
    cpelement_group_441 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(227) & cp_elements(445));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(441),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2004_load_0_req_0 <= cp_elements(441);
    cp_elements(442) <= cp_elements(227);
    ptr_deref_2004_base_resize_req_0 <= cp_elements(442);
    cp_elements(443) <= ptr_deref_2004_base_resize_ack_0;
    ptr_deref_2004_root_address_inst_req_0 <= cp_elements(443);
    cp_elements(444) <= ptr_deref_2004_root_address_inst_ack_0;
    ptr_deref_2004_addr_0_req_0 <= cp_elements(444);
    cp_elements(445) <= ptr_deref_2004_addr_0_ack_0;
    cp_elements(446) <= ptr_deref_2004_load_0_ack_0;
    ptr_deref_2004_load_0_req_1 <= cp_elements(446);
    cp_elements(447) <= ptr_deref_2004_load_0_ack_1;
    ptr_deref_2004_gather_scatter_req_0 <= cp_elements(447);
    cp_elements(448) <= ptr_deref_2004_gather_scatter_ack_0;
    cpelement_group_449 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(448) & cp_elements(450));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(449),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2008_inst_req_0 <= cp_elements(449);
    cp_elements(450) <= cp_elements(206);
    cp_elements(451) <= type_cast_2008_inst_ack_0;
    cpelement_group_452 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(451) & cp_elements(453));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(452),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2014_inst_req_0 <= cp_elements(452);
    cp_elements(453) <= cp_elements(206);
    cp_elements(454) <= binary_2014_inst_ack_0;
    binary_2014_inst_req_1 <= cp_elements(454);
    cp_elements(455) <= binary_2014_inst_ack_1;
    cpelement_group_456 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(350) & cp_elements(365) & cp_elements(457));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(456),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2019_inst_req_0 <= cp_elements(456);
    cp_elements(457) <= cp_elements(206);
    cp_elements(458) <= binary_2019_inst_ack_0;
    binary_2019_inst_req_1 <= cp_elements(458);
    cp_elements(459) <= binary_2019_inst_ack_1;
    cpelement_group_460 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(380) & cp_elements(459) & cp_elements(461));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(460),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2024_inst_req_0 <= cp_elements(460);
    cp_elements(461) <= cp_elements(206);
    cp_elements(462) <= binary_2024_inst_ack_0;
    binary_2024_inst_req_1 <= cp_elements(462);
    cp_elements(463) <= binary_2024_inst_ack_1;
    cpelement_group_464 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(395) & cp_elements(463) & cp_elements(465));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(464),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2029_inst_req_0 <= cp_elements(464);
    cp_elements(465) <= cp_elements(206);
    cp_elements(466) <= binary_2029_inst_ack_0;
    binary_2029_inst_req_1 <= cp_elements(466);
    cp_elements(467) <= binary_2029_inst_ack_1;
    cpelement_group_468 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(410) & cp_elements(467) & cp_elements(469));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(468),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2034_inst_req_0 <= cp_elements(468);
    cp_elements(469) <= cp_elements(206);
    cp_elements(470) <= binary_2034_inst_ack_0;
    binary_2034_inst_req_1 <= cp_elements(470);
    cp_elements(471) <= binary_2034_inst_ack_1;
    cpelement_group_472 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(425) & cp_elements(471) & cp_elements(473));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(472),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2039_inst_req_0 <= cp_elements(472);
    cp_elements(473) <= cp_elements(206);
    cp_elements(474) <= binary_2039_inst_ack_0;
    binary_2039_inst_req_1 <= cp_elements(474);
    cp_elements(475) <= binary_2039_inst_ack_1;
    cpelement_group_476 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(440) & cp_elements(475) & cp_elements(477));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(476),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2044_inst_req_0 <= cp_elements(476);
    cp_elements(477) <= cp_elements(206);
    cp_elements(478) <= binary_2044_inst_ack_0;
    binary_2044_inst_req_1 <= cp_elements(478);
    cp_elements(479) <= binary_2044_inst_ack_1;
    cpelement_group_480 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(455) & cp_elements(479) & cp_elements(481));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(480),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2049_inst_req_0 <= cp_elements(480);
    cp_elements(481) <= cp_elements(206);
    cp_elements(482) <= binary_2049_inst_ack_0;
    binary_2049_inst_req_1 <= cp_elements(482);
    cp_elements(483) <= binary_2049_inst_ack_1;
    cpelement_group_484 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(485) & cp_elements(486));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(484),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2055_inst_req_0 <= cp_elements(484);
    cp_elements(485) <= cp_elements(206);
    cp_elements(486) <= cp_elements(206);
    cp_elements(487) <= binary_2055_inst_ack_0;
    binary_2055_inst_req_1 <= cp_elements(487);
    cp_elements(488) <= binary_2055_inst_ack_1;
    cpelement_group_489 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(483) & cp_elements(488));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(489),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(490) <= cp_elements(2);
    cp_elements(491) <= false;
    cp_elements(492) <= cp_elements(491);
    cp_elements(493) <= cp_elements(2);
    if_stmt_2063_branch_req_0 <= cp_elements(493);
    cp_elements(494) <= cp_elements(493);
    cp_elements(495) <= cp_elements(494);
    cp_elements(496) <= if_stmt_2063_branch_ack_1;
    simple_obj_ref_2091_inst_req_0 <= cp_elements(496);
    cp_elements(497) <= cp_elements(494);
    cp_elements(498) <= if_stmt_2063_branch_ack_0;
    cp_elements(499) <= simple_obj_ref_2070_inst_ack_0;
    simple_obj_ref_2080_inst_req_0 <= cp_elements(499);
    cp_elements(500) <= simple_obj_ref_2080_inst_ack_0;
    cp_elements(501) <= cp_elements(500);
    cpelement_group_502 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(503) & cp_elements(504));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(502),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2087_inst_req_0 <= cp_elements(502);
    cp_elements(503) <= cp_elements(501);
    cp_elements(504) <= cp_elements(501);
    cp_elements(505) <= binary_2087_inst_ack_0;
    binary_2087_inst_req_1 <= cp_elements(505);
    cp_elements(506) <= binary_2087_inst_ack_1;
    type_cast_1819_inst_req_0 <= cp_elements(506);
    cp_elements(507) <= simple_obj_ref_2091_inst_ack_0;
    simple_obj_ref_2101_inst_req_0 <= cp_elements(507);
    cp_elements(508) <= simple_obj_ref_2101_inst_ack_0;
    simple_obj_ref_2110_inst_req_0 <= cp_elements(508);
    cp_elements(509) <= simple_obj_ref_2110_inst_ack_0;
    simple_obj_ref_2120_inst_req_0 <= cp_elements(509);
    cp_elements(510) <= simple_obj_ref_2120_inst_ack_0;
    cp_elements(511) <= OrReduce(cp_elements(0) & cp_elements(510));
    cp_elements(512) <= cp_elements(511);
    simple_obj_ref_1613_inst_req_0 <= cp_elements(512);
    cp_elements(513) <= type_cast_1819_inst_ack_0;
    phi_stmt_1816_req_0 <= cp_elements(513);
    cp_elements(514) <= OrReduce(cp_elements(205) & cp_elements(513));
    cp_elements(515) <= cp_elements(514);
    cp_elements(516) <= phi_stmt_1816_ack_0;
    cp_elements(517) <= false;
    cp_elements(518) <= cp_elements(517);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1622_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1622_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1622_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1635_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1635_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1635_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1654_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1654_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1654_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1673_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1673_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1673_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1692_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1692_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1692_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1711_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1711_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1711_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1744_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1744_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1744_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1838_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1838_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1838_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1838_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1848_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1848_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1848_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1848_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1858_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1858_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1858_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1858_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1868_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1878_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1878_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1878_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1878_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1888_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1898_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1898_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1898_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1898_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1908_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1908_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1908_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1908_root_address : std_logic_vector(10 downto 0);
    signal exitcond_2056 : std_logic_vector(0 downto 0);
    signal iNsTr_10_2100 : std_logic_vector(31 downto 0);
    signal iNsTr_12_2109 : std_logic_vector(31 downto 0);
    signal iNsTr_14_2119 : std_logic_vector(31 downto 0);
    signal iNsTr_18_2079 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1611 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1800 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1810 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2062 : std_logic_vector(31 downto 0);
    signal indvar_1816 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2088 : std_logic_vector(31 downto 0);
    signal ins38_1794 : std_logic_vector(63 downto 0);
    signal ins77_2050 : std_logic_vector(63 downto 0);
    signal mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_1764 : std_logic_vector(63 downto 0);
    signal mask17x_xmaskedx_xmaskedx_xmasked_1769 : std_logic_vector(63 downto 0);
    signal mask22x_xmaskedx_xmaskedx_xmasked_1774 : std_logic_vector(63 downto 0);
    signal mask27x_xmaskedx_xmasked_1779 : std_logic_vector(63 downto 0);
    signal mask32x_xmasked_1784 : std_logic_vector(63 downto 0);
    signal mask37_1789 : std_logic_vector(63 downto 0);
    signal mask51_2020 : std_logic_vector(63 downto 0);
    signal mask56_2025 : std_logic_vector(63 downto 0);
    signal mask61x_xmaskedx_xmasked_2030 : std_logic_vector(63 downto 0);
    signal mask66x_xmaskedx_xmasked_2035 : std_logic_vector(63 downto 0);
    signal mask71x_xmasked_2040 : std_logic_vector(63 downto 0);
    signal mask76_2045 : std_logic_vector(63 downto 0);
    signal ptr_deref_1626_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1626_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1626_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1626_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1626_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1639_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1639_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1639_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1639_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1639_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1658_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1658_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1658_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1658_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1658_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1677_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1677_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1677_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1677_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1677_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1696_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1696_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1696_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1696_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1696_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1715_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1715_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1715_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1715_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1715_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1729_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1729_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1729_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1729_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1729_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1748_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1748_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1748_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1748_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1748_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1912_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1912_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1912_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1912_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1912_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1920_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1920_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1920_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1920_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1920_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1934_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1934_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1934_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1934_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1934_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1948_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1948_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1948_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1948_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1948_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1962_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1962_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1962_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1962_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1962_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1976_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1976_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1976_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1976_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1976_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1990_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1990_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1990_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1990_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1990_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2004_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2004_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2004_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2004_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2004_word_offset_0 : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1837_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1837_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1847_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1847_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1857_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1857_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1867_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1867_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1877_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1877_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1887_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1887_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1897_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1897_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1907_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1907_scaled : std_logic_vector(10 downto 0);
    signal tmp10_1663 : std_logic_vector(63 downto 0);
    signal tmp11_1669 : std_logic_vector(63 downto 0);
    signal tmp124_1618 : std_logic_vector(31 downto 0);
    signal tmp125_1623 : std_logic_vector(31 downto 0);
    signal tmp126_1627 : std_logic_vector(7 downto 0);
    signal tmp127_1636 : std_logic_vector(31 downto 0);
    signal tmp128_1640 : std_logic_vector(7 downto 0);
    signal tmp129_1655 : std_logic_vector(31 downto 0);
    signal tmp130_1659 : std_logic_vector(7 downto 0);
    signal tmp131_1674 : std_logic_vector(31 downto 0);
    signal tmp132_1678 : std_logic_vector(7 downto 0);
    signal tmp133_1693 : std_logic_vector(31 downto 0);
    signal tmp134_1697 : std_logic_vector(7 downto 0);
    signal tmp135_1712 : std_logic_vector(31 downto 0);
    signal tmp136_1716 : std_logic_vector(7 downto 0);
    signal tmp137_1730 : std_logic_vector(7 downto 0);
    signal tmp138_1745 : std_logic_vector(31 downto 0);
    signal tmp139_1749 : std_logic_vector(7 downto 0);
    signal tmp146_1909 : std_logic_vector(31 downto 0);
    signal tmp147_1913 : std_logic_vector(7 downto 0);
    signal tmp151_1899 : std_logic_vector(31 downto 0);
    signal tmp152_1921 : std_logic_vector(7 downto 0);
    signal tmp156_1889 : std_logic_vector(31 downto 0);
    signal tmp157_1935 : std_logic_vector(7 downto 0);
    signal tmp15_1682 : std_logic_vector(63 downto 0);
    signal tmp161_1879 : std_logic_vector(31 downto 0);
    signal tmp162_1949 : std_logic_vector(7 downto 0);
    signal tmp166_1869 : std_logic_vector(31 downto 0);
    signal tmp167_1963 : std_logic_vector(7 downto 0);
    signal tmp16_1688 : std_logic_vector(63 downto 0);
    signal tmp171_1859 : std_logic_vector(31 downto 0);
    signal tmp172_1977 : std_logic_vector(7 downto 0);
    signal tmp176_1849 : std_logic_vector(31 downto 0);
    signal tmp177_1991 : std_logic_vector(7 downto 0);
    signal tmp180_1839 : std_logic_vector(31 downto 0);
    signal tmp181_2005 : std_logic_vector(7 downto 0);
    signal tmp20_1701 : std_logic_vector(63 downto 0);
    signal tmp21_1707 : std_logic_vector(63 downto 0);
    signal tmp224_1829 : std_logic_vector(31 downto 0);
    signal tmp225_1835 : std_logic_vector(31 downto 0);
    signal tmp226_1845 : std_logic_vector(31 downto 0);
    signal tmp227_1855 : std_logic_vector(31 downto 0);
    signal tmp228_1865 : std_logic_vector(31 downto 0);
    signal tmp229_1875 : std_logic_vector(31 downto 0);
    signal tmp230_1885 : std_logic_vector(31 downto 0);
    signal tmp231_1895 : std_logic_vector(31 downto 0);
    signal tmp232_1905 : std_logic_vector(31 downto 0);
    signal tmp25_1720 : std_logic_vector(63 downto 0);
    signal tmp26_1726 : std_logic_vector(63 downto 0);
    signal tmp30_1734 : std_logic_vector(63 downto 0);
    signal tmp31_1740 : std_logic_vector(63 downto 0);
    signal tmp35_1753 : std_logic_vector(63 downto 0);
    signal tmp36_1759 : std_logic_vector(63 downto 0);
    signal tmp3_1631 : std_logic_vector(63 downto 0);
    signal tmp40_1917 : std_logic_vector(63 downto 0);
    signal tmp44_1925 : std_logic_vector(63 downto 0);
    signal tmp45_1931 : std_logic_vector(63 downto 0);
    signal tmp49_1939 : std_logic_vector(63 downto 0);
    signal tmp50_1945 : std_logic_vector(63 downto 0);
    signal tmp54_1953 : std_logic_vector(63 downto 0);
    signal tmp55_1959 : std_logic_vector(63 downto 0);
    signal tmp59_1967 : std_logic_vector(63 downto 0);
    signal tmp5_1644 : std_logic_vector(63 downto 0);
    signal tmp60_1973 : std_logic_vector(63 downto 0);
    signal tmp64_1981 : std_logic_vector(63 downto 0);
    signal tmp65_1987 : std_logic_vector(63 downto 0);
    signal tmp69_1995 : std_logic_vector(63 downto 0);
    signal tmp6_1650 : std_logic_vector(63 downto 0);
    signal tmp70_2001 : std_logic_vector(63 downto 0);
    signal tmp74_2009 : std_logic_vector(63 downto 0);
    signal tmp75_2015 : std_logic_vector(63 downto 0);
    signal tmp_1614 : std_logic_vector(31 downto 0);
    signal type_cast_1648_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1667_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1686_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1705_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1724_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1738_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1757_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1803_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1819_wire : std_logic_vector(31 downto 0);
    signal type_cast_1822_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1827_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1843_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1853_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1863_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1873_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1883_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1893_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1903_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1929_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1957_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1971_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1985_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1999_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2013_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2054_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2072_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2086_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2093_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2112_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1622_final_offset <= "00000000111";
    array_obj_ref_1635_final_offset <= "00000000110";
    array_obj_ref_1654_final_offset <= "00000000101";
    array_obj_ref_1673_final_offset <= "00000000100";
    array_obj_ref_1692_final_offset <= "00000000011";
    array_obj_ref_1711_final_offset <= "00000000010";
    array_obj_ref_1744_final_offset <= "00000000001";
    array_obj_ref_1838_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1848_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1858_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1868_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1878_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1888_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1898_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1908_offset_scale_factor_0 <= "00000000001";
    iNsTr_10_2100 <= "00000000000000000000000000000000";
    iNsTr_12_2109 <= "00000000000000000000000000000000";
    iNsTr_14_2119 <= "00000000000000000000000000000000";
    iNsTr_18_2079 <= "00000000000000000000000000000000";
    iNsTr_1_1611 <= "00000000000000000000000000000000";
    iNsTr_2_1800 <= "00000000000000000000000000000000";
    iNsTr_4_1810 <= "00000000000000000000000000000000";
    iNsTr_7_2062 <= "00000000000000000000000000000000";
    ptr_deref_1626_word_offset_0 <= "00000000000";
    ptr_deref_1639_word_offset_0 <= "00000000000";
    ptr_deref_1658_word_offset_0 <= "00000000000";
    ptr_deref_1677_word_offset_0 <= "00000000000";
    ptr_deref_1696_word_offset_0 <= "00000000000";
    ptr_deref_1715_word_offset_0 <= "00000000000";
    ptr_deref_1729_word_offset_0 <= "00000000000";
    ptr_deref_1748_word_offset_0 <= "00000000000";
    ptr_deref_1912_word_offset_0 <= "00000000000";
    ptr_deref_1920_word_offset_0 <= "00000000000";
    ptr_deref_1934_word_offset_0 <= "00000000000";
    ptr_deref_1948_word_offset_0 <= "00000000000";
    ptr_deref_1962_word_offset_0 <= "00000000000";
    ptr_deref_1976_word_offset_0 <= "00000000000";
    ptr_deref_1990_word_offset_0 <= "00000000000";
    ptr_deref_2004_word_offset_0 <= "00000000000";
    type_cast_1648_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1667_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1686_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1705_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1738_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1757_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1803_wire_constant <= "11111111";
    type_cast_1822_wire_constant <= "00000000000000000000000000000000";
    type_cast_1827_wire_constant <= "00000000000000000000000000000011";
    type_cast_1833_wire_constant <= "00000000000000000000000000001000";
    type_cast_1843_wire_constant <= "00000000000000000000000000001001";
    type_cast_1853_wire_constant <= "00000000000000000000000000001010";
    type_cast_1863_wire_constant <= "00000000000000000000000000001011";
    type_cast_1873_wire_constant <= "00000000000000000000000000001100";
    type_cast_1883_wire_constant <= "00000000000000000000000000001101";
    type_cast_1893_wire_constant <= "00000000000000000000000000001110";
    type_cast_1903_wire_constant <= "00000000000000000000000000001111";
    type_cast_1929_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1957_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1971_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1985_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1999_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2013_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2054_wire_constant <= "00000000000000000000000000011110";
    type_cast_2072_wire_constant <= "00000000";
    type_cast_2086_wire_constant <= "00000000000000000000000000000001";
    type_cast_2093_wire_constant <= "00000001";
    type_cast_2112_wire_constant <= "00000001";
    phi_stmt_1816: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1819_wire & type_cast_1822_wire_constant;
      req <= phi_stmt_1816_req_0 & phi_stmt_1816_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1816_ack_0,
          idata => idata,
          odata => indvar_1816,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1816
    array_obj_ref_1622_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1622_resized_base_address, req => array_obj_ref_1622_base_resize_req_0, ack => array_obj_ref_1622_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1622_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1622_root_address, dout => tmp125_1623, req => array_obj_ref_1622_final_reg_req_0, ack => array_obj_ref_1622_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1635_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1635_resized_base_address, req => array_obj_ref_1635_base_resize_req_0, ack => array_obj_ref_1635_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1635_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1635_root_address, dout => tmp127_1636, req => array_obj_ref_1635_final_reg_req_0, ack => array_obj_ref_1635_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1654_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1654_resized_base_address, req => array_obj_ref_1654_base_resize_req_0, ack => array_obj_ref_1654_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1654_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1654_root_address, dout => tmp129_1655, req => array_obj_ref_1654_final_reg_req_0, ack => array_obj_ref_1654_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1673_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1673_resized_base_address, req => array_obj_ref_1673_base_resize_req_0, ack => array_obj_ref_1673_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1673_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1673_root_address, dout => tmp131_1674, req => array_obj_ref_1673_final_reg_req_0, ack => array_obj_ref_1673_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1692_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1692_resized_base_address, req => array_obj_ref_1692_base_resize_req_0, ack => array_obj_ref_1692_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1692_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1692_root_address, dout => tmp133_1693, req => array_obj_ref_1692_final_reg_req_0, ack => array_obj_ref_1692_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1711_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1711_resized_base_address, req => array_obj_ref_1711_base_resize_req_0, ack => array_obj_ref_1711_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1711_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1711_root_address, dout => tmp135_1712, req => array_obj_ref_1711_final_reg_req_0, ack => array_obj_ref_1711_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1744_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1744_resized_base_address, req => array_obj_ref_1744_base_resize_req_0, ack => array_obj_ref_1744_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1744_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1744_root_address, dout => tmp138_1745, req => array_obj_ref_1744_final_reg_req_0, ack => array_obj_ref_1744_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1838_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1838_resized_base_address, req => array_obj_ref_1838_base_resize_req_0, ack => array_obj_ref_1838_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1838_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1838_root_address, dout => tmp180_1839, req => array_obj_ref_1838_final_reg_req_0, ack => array_obj_ref_1838_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1838_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp225_1835, dout => simple_obj_ref_1837_resized, req => array_obj_ref_1838_index_0_resize_req_0, ack => array_obj_ref_1838_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1838_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1837_scaled, dout => array_obj_ref_1838_final_offset, req => array_obj_ref_1838_offset_inst_req_0, ack => array_obj_ref_1838_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1848_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1848_resized_base_address, req => array_obj_ref_1848_base_resize_req_0, ack => array_obj_ref_1848_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1848_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1848_root_address, dout => tmp176_1849, req => array_obj_ref_1848_final_reg_req_0, ack => array_obj_ref_1848_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1848_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp226_1845, dout => simple_obj_ref_1847_resized, req => array_obj_ref_1848_index_0_resize_req_0, ack => array_obj_ref_1848_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1848_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1847_scaled, dout => array_obj_ref_1848_final_offset, req => array_obj_ref_1848_offset_inst_req_0, ack => array_obj_ref_1848_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1858_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1858_resized_base_address, req => array_obj_ref_1858_base_resize_req_0, ack => array_obj_ref_1858_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1858_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1858_root_address, dout => tmp171_1859, req => array_obj_ref_1858_final_reg_req_0, ack => array_obj_ref_1858_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1858_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp227_1855, dout => simple_obj_ref_1857_resized, req => array_obj_ref_1858_index_0_resize_req_0, ack => array_obj_ref_1858_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1858_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1857_scaled, dout => array_obj_ref_1858_final_offset, req => array_obj_ref_1858_offset_inst_req_0, ack => array_obj_ref_1858_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1868_resized_base_address, req => array_obj_ref_1868_base_resize_req_0, ack => array_obj_ref_1868_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1868_root_address, dout => tmp166_1869, req => array_obj_ref_1868_final_reg_req_0, ack => array_obj_ref_1868_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp228_1865, dout => simple_obj_ref_1867_resized, req => array_obj_ref_1868_index_0_resize_req_0, ack => array_obj_ref_1868_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1868_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1867_scaled, dout => array_obj_ref_1868_final_offset, req => array_obj_ref_1868_offset_inst_req_0, ack => array_obj_ref_1868_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1878_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1878_resized_base_address, req => array_obj_ref_1878_base_resize_req_0, ack => array_obj_ref_1878_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1878_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1878_root_address, dout => tmp161_1879, req => array_obj_ref_1878_final_reg_req_0, ack => array_obj_ref_1878_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1878_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp229_1875, dout => simple_obj_ref_1877_resized, req => array_obj_ref_1878_index_0_resize_req_0, ack => array_obj_ref_1878_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1878_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1877_scaled, dout => array_obj_ref_1878_final_offset, req => array_obj_ref_1878_offset_inst_req_0, ack => array_obj_ref_1878_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1888_resized_base_address, req => array_obj_ref_1888_base_resize_req_0, ack => array_obj_ref_1888_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1888_root_address, dout => tmp156_1889, req => array_obj_ref_1888_final_reg_req_0, ack => array_obj_ref_1888_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp230_1885, dout => simple_obj_ref_1887_resized, req => array_obj_ref_1888_index_0_resize_req_0, ack => array_obj_ref_1888_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1887_scaled, dout => array_obj_ref_1888_final_offset, req => array_obj_ref_1888_offset_inst_req_0, ack => array_obj_ref_1888_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1898_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1898_resized_base_address, req => array_obj_ref_1898_base_resize_req_0, ack => array_obj_ref_1898_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1898_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1898_root_address, dout => tmp151_1899, req => array_obj_ref_1898_final_reg_req_0, ack => array_obj_ref_1898_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1898_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp231_1895, dout => simple_obj_ref_1897_resized, req => array_obj_ref_1898_index_0_resize_req_0, ack => array_obj_ref_1898_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1898_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1897_scaled, dout => array_obj_ref_1898_final_offset, req => array_obj_ref_1898_offset_inst_req_0, ack => array_obj_ref_1898_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1908_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => array_obj_ref_1908_resized_base_address, req => array_obj_ref_1908_base_resize_req_0, ack => array_obj_ref_1908_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1908_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1908_root_address, dout => tmp146_1909, req => array_obj_ref_1908_final_reg_req_0, ack => array_obj_ref_1908_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1908_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp232_1905, dout => simple_obj_ref_1907_resized, req => array_obj_ref_1908_index_0_resize_req_0, ack => array_obj_ref_1908_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1908_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1907_scaled, dout => array_obj_ref_1908_final_offset, req => array_obj_ref_1908_offset_inst_req_0, ack => array_obj_ref_1908_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1626_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp125_1623, dout => ptr_deref_1626_resized_base_address, req => ptr_deref_1626_base_resize_req_0, ack => ptr_deref_1626_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1639_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp127_1636, dout => ptr_deref_1639_resized_base_address, req => ptr_deref_1639_base_resize_req_0, ack => ptr_deref_1639_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1658_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp129_1655, dout => ptr_deref_1658_resized_base_address, req => ptr_deref_1658_base_resize_req_0, ack => ptr_deref_1658_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1677_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp131_1674, dout => ptr_deref_1677_resized_base_address, req => ptr_deref_1677_base_resize_req_0, ack => ptr_deref_1677_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1696_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp133_1693, dout => ptr_deref_1696_resized_base_address, req => ptr_deref_1696_base_resize_req_0, ack => ptr_deref_1696_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1715_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp135_1712, dout => ptr_deref_1715_resized_base_address, req => ptr_deref_1715_base_resize_req_0, ack => ptr_deref_1715_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1729_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1618, dout => ptr_deref_1729_resized_base_address, req => ptr_deref_1729_base_resize_req_0, ack => ptr_deref_1729_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1748_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp138_1745, dout => ptr_deref_1748_resized_base_address, req => ptr_deref_1748_base_resize_req_0, ack => ptr_deref_1748_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1912_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp146_1909, dout => ptr_deref_1912_resized_base_address, req => ptr_deref_1912_base_resize_req_0, ack => ptr_deref_1912_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1920_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp151_1899, dout => ptr_deref_1920_resized_base_address, req => ptr_deref_1920_base_resize_req_0, ack => ptr_deref_1920_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1934_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp156_1889, dout => ptr_deref_1934_resized_base_address, req => ptr_deref_1934_base_resize_req_0, ack => ptr_deref_1934_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1948_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp161_1879, dout => ptr_deref_1948_resized_base_address, req => ptr_deref_1948_base_resize_req_0, ack => ptr_deref_1948_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1962_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp166_1869, dout => ptr_deref_1962_resized_base_address, req => ptr_deref_1962_base_resize_req_0, ack => ptr_deref_1962_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1976_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp171_1859, dout => ptr_deref_1976_resized_base_address, req => ptr_deref_1976_base_resize_req_0, ack => ptr_deref_1976_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1990_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp176_1849, dout => ptr_deref_1990_resized_base_address, req => ptr_deref_1990_base_resize_req_0, ack => ptr_deref_1990_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2004_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp180_1839, dout => ptr_deref_2004_resized_base_address, req => ptr_deref_2004_base_resize_req_0, ack => ptr_deref_2004_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1617_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_1614, dout => tmp124_1618, req => type_cast_1617_inst_req_0, ack => type_cast_1617_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1630_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp126_1627, dout => tmp3_1631, req => type_cast_1630_inst_req_0, ack => type_cast_1630_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1643_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp128_1640, dout => tmp5_1644, req => type_cast_1643_inst_req_0, ack => type_cast_1643_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1662_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp130_1659, dout => tmp10_1663, req => type_cast_1662_inst_req_0, ack => type_cast_1662_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1681_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp132_1678, dout => tmp15_1682, req => type_cast_1681_inst_req_0, ack => type_cast_1681_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1700_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp134_1697, dout => tmp20_1701, req => type_cast_1700_inst_req_0, ack => type_cast_1700_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1719_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp136_1716, dout => tmp25_1720, req => type_cast_1719_inst_req_0, ack => type_cast_1719_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1733_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp137_1730, dout => tmp30_1734, req => type_cast_1733_inst_req_0, ack => type_cast_1733_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1752_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp139_1749, dout => tmp35_1753, req => type_cast_1752_inst_req_0, ack => type_cast_1752_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1819_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => indvarx_xnext_2088, dout => type_cast_1819_wire, req => type_cast_1819_inst_req_0, ack => type_cast_1819_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1916_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp147_1913, dout => tmp40_1917, req => type_cast_1916_inst_req_0, ack => type_cast_1916_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1924_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp152_1921, dout => tmp44_1925, req => type_cast_1924_inst_req_0, ack => type_cast_1924_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1938_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp157_1935, dout => tmp49_1939, req => type_cast_1938_inst_req_0, ack => type_cast_1938_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1952_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp162_1949, dout => tmp54_1953, req => type_cast_1952_inst_req_0, ack => type_cast_1952_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1966_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp167_1963, dout => tmp59_1967, req => type_cast_1966_inst_req_0, ack => type_cast_1966_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1980_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp172_1977, dout => tmp64_1981, req => type_cast_1980_inst_req_0, ack => type_cast_1980_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1994_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp177_1991, dout => tmp69_1995, req => type_cast_1994_inst_req_0, ack => type_cast_1994_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2008_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp181_2005, dout => tmp74_2009, req => type_cast_2008_inst_req_0, ack => type_cast_2008_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1838_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1838_index_0_rename_ack_0 <= array_obj_ref_1838_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1837_resized;
      simple_obj_ref_1837_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1848_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1848_index_0_rename_ack_0 <= array_obj_ref_1848_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1847_resized;
      simple_obj_ref_1847_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1858_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1858_index_0_rename_ack_0 <= array_obj_ref_1858_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1857_resized;
      simple_obj_ref_1857_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1868_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1868_index_0_rename_ack_0 <= array_obj_ref_1868_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1867_resized;
      simple_obj_ref_1867_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1878_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1878_index_0_rename_ack_0 <= array_obj_ref_1878_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1877_resized;
      simple_obj_ref_1877_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1888_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1888_index_0_rename_ack_0 <= array_obj_ref_1888_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1887_resized;
      simple_obj_ref_1887_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1898_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1898_index_0_rename_ack_0 <= array_obj_ref_1898_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1897_resized;
      simple_obj_ref_1897_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1908_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1908_index_0_rename_ack_0 <= array_obj_ref_1908_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1907_resized;
      simple_obj_ref_1907_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1626_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1626_addr_0_ack_0 <= ptr_deref_1626_addr_0_req_0;
      aggregated_sig <= ptr_deref_1626_root_address;
      ptr_deref_1626_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1626_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1626_gather_scatter_ack_0 <= ptr_deref_1626_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1626_data_0;
      tmp126_1627 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1626_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1626_root_address_inst_ack_0 <= ptr_deref_1626_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1626_resized_base_address;
      ptr_deref_1626_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1639_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1639_addr_0_ack_0 <= ptr_deref_1639_addr_0_req_0;
      aggregated_sig <= ptr_deref_1639_root_address;
      ptr_deref_1639_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1639_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1639_gather_scatter_ack_0 <= ptr_deref_1639_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1639_data_0;
      tmp128_1640 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1639_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1639_root_address_inst_ack_0 <= ptr_deref_1639_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1639_resized_base_address;
      ptr_deref_1639_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1658_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1658_addr_0_ack_0 <= ptr_deref_1658_addr_0_req_0;
      aggregated_sig <= ptr_deref_1658_root_address;
      ptr_deref_1658_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1658_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1658_gather_scatter_ack_0 <= ptr_deref_1658_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1658_data_0;
      tmp130_1659 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1658_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1658_root_address_inst_ack_0 <= ptr_deref_1658_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1658_resized_base_address;
      ptr_deref_1658_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1677_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1677_addr_0_ack_0 <= ptr_deref_1677_addr_0_req_0;
      aggregated_sig <= ptr_deref_1677_root_address;
      ptr_deref_1677_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1677_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1677_gather_scatter_ack_0 <= ptr_deref_1677_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1677_data_0;
      tmp132_1678 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1677_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1677_root_address_inst_ack_0 <= ptr_deref_1677_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1677_resized_base_address;
      ptr_deref_1677_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1696_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1696_addr_0_ack_0 <= ptr_deref_1696_addr_0_req_0;
      aggregated_sig <= ptr_deref_1696_root_address;
      ptr_deref_1696_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1696_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1696_gather_scatter_ack_0 <= ptr_deref_1696_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1696_data_0;
      tmp134_1697 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1696_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1696_root_address_inst_ack_0 <= ptr_deref_1696_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1696_resized_base_address;
      ptr_deref_1696_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1715_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1715_addr_0_ack_0 <= ptr_deref_1715_addr_0_req_0;
      aggregated_sig <= ptr_deref_1715_root_address;
      ptr_deref_1715_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1715_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1715_gather_scatter_ack_0 <= ptr_deref_1715_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1715_data_0;
      tmp136_1716 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1715_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1715_root_address_inst_ack_0 <= ptr_deref_1715_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1715_resized_base_address;
      ptr_deref_1715_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1729_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1729_addr_0_ack_0 <= ptr_deref_1729_addr_0_req_0;
      aggregated_sig <= ptr_deref_1729_root_address;
      ptr_deref_1729_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1729_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1729_gather_scatter_ack_0 <= ptr_deref_1729_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1729_data_0;
      tmp137_1730 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1729_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1729_root_address_inst_ack_0 <= ptr_deref_1729_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1729_resized_base_address;
      ptr_deref_1729_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1748_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1748_addr_0_ack_0 <= ptr_deref_1748_addr_0_req_0;
      aggregated_sig <= ptr_deref_1748_root_address;
      ptr_deref_1748_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1748_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1748_gather_scatter_ack_0 <= ptr_deref_1748_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1748_data_0;
      tmp139_1749 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1748_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1748_root_address_inst_ack_0 <= ptr_deref_1748_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1748_resized_base_address;
      ptr_deref_1748_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1912_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1912_addr_0_ack_0 <= ptr_deref_1912_addr_0_req_0;
      aggregated_sig <= ptr_deref_1912_root_address;
      ptr_deref_1912_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1912_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1912_gather_scatter_ack_0 <= ptr_deref_1912_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1912_data_0;
      tmp147_1913 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1912_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1912_root_address_inst_ack_0 <= ptr_deref_1912_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1912_resized_base_address;
      ptr_deref_1912_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1920_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1920_addr_0_ack_0 <= ptr_deref_1920_addr_0_req_0;
      aggregated_sig <= ptr_deref_1920_root_address;
      ptr_deref_1920_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1920_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1920_gather_scatter_ack_0 <= ptr_deref_1920_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1920_data_0;
      tmp152_1921 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1920_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1920_root_address_inst_ack_0 <= ptr_deref_1920_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1920_resized_base_address;
      ptr_deref_1920_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1934_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1934_addr_0_ack_0 <= ptr_deref_1934_addr_0_req_0;
      aggregated_sig <= ptr_deref_1934_root_address;
      ptr_deref_1934_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1934_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1934_gather_scatter_ack_0 <= ptr_deref_1934_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1934_data_0;
      tmp157_1935 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1934_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1934_root_address_inst_ack_0 <= ptr_deref_1934_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1934_resized_base_address;
      ptr_deref_1934_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1948_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1948_addr_0_ack_0 <= ptr_deref_1948_addr_0_req_0;
      aggregated_sig <= ptr_deref_1948_root_address;
      ptr_deref_1948_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1948_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1948_gather_scatter_ack_0 <= ptr_deref_1948_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1948_data_0;
      tmp162_1949 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1948_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1948_root_address_inst_ack_0 <= ptr_deref_1948_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1948_resized_base_address;
      ptr_deref_1948_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1962_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1962_addr_0_ack_0 <= ptr_deref_1962_addr_0_req_0;
      aggregated_sig <= ptr_deref_1962_root_address;
      ptr_deref_1962_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1962_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1962_gather_scatter_ack_0 <= ptr_deref_1962_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1962_data_0;
      tmp167_1963 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1962_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1962_root_address_inst_ack_0 <= ptr_deref_1962_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1962_resized_base_address;
      ptr_deref_1962_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1976_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1976_addr_0_ack_0 <= ptr_deref_1976_addr_0_req_0;
      aggregated_sig <= ptr_deref_1976_root_address;
      ptr_deref_1976_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1976_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1976_gather_scatter_ack_0 <= ptr_deref_1976_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1976_data_0;
      tmp172_1977 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1976_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1976_root_address_inst_ack_0 <= ptr_deref_1976_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1976_resized_base_address;
      ptr_deref_1976_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1990_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1990_addr_0_ack_0 <= ptr_deref_1990_addr_0_req_0;
      aggregated_sig <= ptr_deref_1990_root_address;
      ptr_deref_1990_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1990_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1990_gather_scatter_ack_0 <= ptr_deref_1990_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1990_data_0;
      tmp177_1991 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1990_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1990_root_address_inst_ack_0 <= ptr_deref_1990_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1990_resized_base_address;
      ptr_deref_1990_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2004_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2004_addr_0_ack_0 <= ptr_deref_2004_addr_0_req_0;
      aggregated_sig <= ptr_deref_2004_root_address;
      ptr_deref_2004_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2004_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2004_gather_scatter_ack_0 <= ptr_deref_2004_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2004_data_0;
      tmp181_2005 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2004_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2004_root_address_inst_ack_0 <= ptr_deref_2004_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2004_resized_base_address;
      ptr_deref_2004_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    if_stmt_2063_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_2056;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2063_branch_req_0,
          ack0 => if_stmt_2063_branch_ack_0,
          ack1 => if_stmt_2063_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1622_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1622_resized_base_address;
      array_obj_ref_1622_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000111",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1622_root_address_inst_req_0,
          ackL => array_obj_ref_1622_root_address_inst_ack_0,
          reqR => array_obj_ref_1622_root_address_inst_req_1,
          ackR => array_obj_ref_1622_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1635_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1635_resized_base_address;
      array_obj_ref_1635_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000110",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1635_root_address_inst_req_0,
          ackL => array_obj_ref_1635_root_address_inst_ack_0,
          reqR => array_obj_ref_1635_root_address_inst_req_1,
          ackR => array_obj_ref_1635_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1654_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1654_resized_base_address;
      array_obj_ref_1654_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000101",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1654_root_address_inst_req_0,
          ackL => array_obj_ref_1654_root_address_inst_ack_0,
          reqR => array_obj_ref_1654_root_address_inst_req_1,
          ackR => array_obj_ref_1654_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1673_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1673_resized_base_address;
      array_obj_ref_1673_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1673_root_address_inst_req_0,
          ackL => array_obj_ref_1673_root_address_inst_ack_0,
          reqR => array_obj_ref_1673_root_address_inst_req_1,
          ackR => array_obj_ref_1673_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1692_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1692_resized_base_address;
      array_obj_ref_1692_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000011",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1692_root_address_inst_req_0,
          ackL => array_obj_ref_1692_root_address_inst_ack_0,
          reqR => array_obj_ref_1692_root_address_inst_req_1,
          ackR => array_obj_ref_1692_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1711_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1711_resized_base_address;
      array_obj_ref_1711_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000010",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1711_root_address_inst_req_0,
          ackL => array_obj_ref_1711_root_address_inst_ack_0,
          reqR => array_obj_ref_1711_root_address_inst_req_1,
          ackR => array_obj_ref_1711_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1744_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1744_resized_base_address;
      array_obj_ref_1744_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1744_root_address_inst_req_0,
          ackL => array_obj_ref_1744_root_address_inst_ack_0,
          reqR => array_obj_ref_1744_root_address_inst_req_1,
          ackR => array_obj_ref_1744_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_1838_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1838_final_offset & array_obj_ref_1838_resized_base_address;
      array_obj_ref_1838_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1838_root_address_inst_req_0,
          ackL => array_obj_ref_1838_root_address_inst_ack_0,
          reqR => array_obj_ref_1838_root_address_inst_req_1,
          ackR => array_obj_ref_1838_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_1848_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1848_final_offset & array_obj_ref_1848_resized_base_address;
      array_obj_ref_1848_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1848_root_address_inst_req_0,
          ackL => array_obj_ref_1848_root_address_inst_ack_0,
          reqR => array_obj_ref_1848_root_address_inst_req_1,
          ackR => array_obj_ref_1848_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_1858_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1858_final_offset & array_obj_ref_1858_resized_base_address;
      array_obj_ref_1858_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1858_root_address_inst_req_0,
          ackL => array_obj_ref_1858_root_address_inst_ack_0,
          reqR => array_obj_ref_1858_root_address_inst_req_1,
          ackR => array_obj_ref_1858_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_1868_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1868_final_offset & array_obj_ref_1868_resized_base_address;
      array_obj_ref_1868_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1868_root_address_inst_req_0,
          ackL => array_obj_ref_1868_root_address_inst_ack_0,
          reqR => array_obj_ref_1868_root_address_inst_req_1,
          ackR => array_obj_ref_1868_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_1878_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1878_final_offset & array_obj_ref_1878_resized_base_address;
      array_obj_ref_1878_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1878_root_address_inst_req_0,
          ackL => array_obj_ref_1878_root_address_inst_ack_0,
          reqR => array_obj_ref_1878_root_address_inst_req_1,
          ackR => array_obj_ref_1878_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_1888_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1888_final_offset & array_obj_ref_1888_resized_base_address;
      array_obj_ref_1888_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1888_root_address_inst_req_0,
          ackL => array_obj_ref_1888_root_address_inst_ack_0,
          reqR => array_obj_ref_1888_root_address_inst_req_1,
          ackR => array_obj_ref_1888_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_1898_root_address_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1898_final_offset & array_obj_ref_1898_resized_base_address;
      array_obj_ref_1898_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1898_root_address_inst_req_0,
          ackL => array_obj_ref_1898_root_address_inst_ack_0,
          reqR => array_obj_ref_1898_root_address_inst_req_1,
          ackR => array_obj_ref_1898_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_1908_root_address_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1908_final_offset & array_obj_ref_1908_resized_base_address;
      array_obj_ref_1908_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1908_root_address_inst_req_0,
          ackL => array_obj_ref_1908_root_address_inst_ack_0,
          reqR => array_obj_ref_1908_root_address_inst_req_1,
          ackR => array_obj_ref_1908_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1649_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp5_1644;
      tmp6_1650 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1649_inst_req_0,
          ackL => binary_1649_inst_ack_0,
          reqR => binary_1649_inst_req_1,
          ackR => binary_1649_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1668_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp10_1663;
      tmp11_1669 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1668_inst_req_0,
          ackL => binary_1668_inst_ack_0,
          reqR => binary_1668_inst_req_1,
          ackR => binary_1668_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1687_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_1682;
      tmp16_1688 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1687_inst_req_0,
          ackL => binary_1687_inst_ack_0,
          reqR => binary_1687_inst_req_1,
          ackR => binary_1687_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_1706_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_1701;
      tmp21_1707 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1706_inst_req_0,
          ackL => binary_1706_inst_ack_0,
          reqR => binary_1706_inst_req_1,
          ackR => binary_1706_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_1725_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp25_1720;
      tmp26_1726 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1725_inst_req_0,
          ackL => binary_1725_inst_ack_0,
          reqR => binary_1725_inst_req_1,
          ackR => binary_1725_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_1739_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_1734;
      tmp31_1740 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1739_inst_req_0,
          ackL => binary_1739_inst_ack_0,
          reqR => binary_1739_inst_req_1,
          ackR => binary_1739_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1758_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp35_1753;
      tmp36_1759 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1758_inst_req_0,
          ackL => binary_1758_inst_ack_0,
          reqR => binary_1758_inst_req_1,
          ackR => binary_1758_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1763_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_1650 & tmp3_1631;
      mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_1764 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1763_inst_req_0,
          ackL => binary_1763_inst_ack_0,
          reqR => binary_1763_inst_req_1,
          ackR => binary_1763_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1768_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_1764 & tmp11_1669;
      mask17x_xmaskedx_xmaskedx_xmasked_1769 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1768_inst_req_0,
          ackL => binary_1768_inst_ack_0,
          reqR => binary_1768_inst_req_1,
          ackR => binary_1768_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1773_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask17x_xmaskedx_xmaskedx_xmasked_1769 & tmp16_1688;
      mask22x_xmaskedx_xmaskedx_xmasked_1774 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1773_inst_req_0,
          ackL => binary_1773_inst_ack_0,
          reqR => binary_1773_inst_req_1,
          ackR => binary_1773_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1778_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask22x_xmaskedx_xmaskedx_xmasked_1774 & tmp21_1707;
      mask27x_xmaskedx_xmasked_1779 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1778_inst_req_0,
          ackL => binary_1778_inst_ack_0,
          reqR => binary_1778_inst_req_1,
          ackR => binary_1778_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1783_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask27x_xmaskedx_xmasked_1779 & tmp26_1726;
      mask32x_xmasked_1784 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1783_inst_req_0,
          ackL => binary_1783_inst_ack_0,
          reqR => binary_1783_inst_req_1,
          ackR => binary_1783_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_1788_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask32x_xmasked_1784 & tmp31_1740;
      mask37_1789 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1788_inst_req_0,
          ackL => binary_1788_inst_ack_0,
          reqR => binary_1788_inst_req_1,
          ackR => binary_1788_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_1793_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask37_1789 & tmp36_1759;
      ins38_1794 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1793_inst_req_0,
          ackL => binary_1793_inst_ack_0,
          reqR => binary_1793_inst_req_1,
          ackR => binary_1793_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_1828_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_1816;
      tmp224_1829 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1828_inst_req_0,
          ackL => binary_1828_inst_ack_0,
          reqR => binary_1828_inst_req_1,
          ackR => binary_1828_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_1834_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp225_1835 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1834_inst_req_0,
          ackL => binary_1834_inst_ack_0,
          reqR => binary_1834_inst_req_1,
          ackR => binary_1834_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_1844_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp226_1845 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1844_inst_req_0,
          ackL => binary_1844_inst_ack_0,
          reqR => binary_1844_inst_req_1,
          ackR => binary_1844_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_1854_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp227_1855 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1854_inst_req_0,
          ackL => binary_1854_inst_ack_0,
          reqR => binary_1854_inst_req_1,
          ackR => binary_1854_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_1864_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp228_1865 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1864_inst_req_0,
          ackL => binary_1864_inst_ack_0,
          reqR => binary_1864_inst_req_1,
          ackR => binary_1864_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_1874_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp229_1875 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1874_inst_req_0,
          ackL => binary_1874_inst_ack_0,
          reqR => binary_1874_inst_req_1,
          ackR => binary_1874_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_1884_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp230_1885 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1884_inst_req_0,
          ackL => binary_1884_inst_ack_0,
          reqR => binary_1884_inst_req_1,
          ackR => binary_1884_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_1894_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp231_1895 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1894_inst_req_0,
          ackL => binary_1894_inst_ack_0,
          reqR => binary_1894_inst_req_1,
          ackR => binary_1894_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_1904_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp224_1829;
      tmp232_1905 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1904_inst_req_0,
          ackL => binary_1904_inst_ack_0,
          reqR => binary_1904_inst_req_1,
          ackR => binary_1904_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_1930_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp44_1925;
      tmp45_1931 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1930_inst_req_0,
          ackL => binary_1930_inst_ack_0,
          reqR => binary_1930_inst_req_1,
          ackR => binary_1930_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_1944_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp49_1939;
      tmp50_1945 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1944_inst_req_0,
          ackL => binary_1944_inst_ack_0,
          reqR => binary_1944_inst_req_1,
          ackR => binary_1944_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_1958_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp54_1953;
      tmp55_1959 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1958_inst_req_0,
          ackL => binary_1958_inst_ack_0,
          reqR => binary_1958_inst_req_1,
          ackR => binary_1958_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_1972_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp59_1967;
      tmp60_1973 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1972_inst_req_0,
          ackL => binary_1972_inst_ack_0,
          reqR => binary_1972_inst_req_1,
          ackR => binary_1972_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_1986_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp64_1981;
      tmp65_1987 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1986_inst_req_0,
          ackL => binary_1986_inst_ack_0,
          reqR => binary_1986_inst_req_1,
          ackR => binary_1986_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_2000_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp69_1995;
      tmp70_2001 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2000_inst_req_0,
          ackL => binary_2000_inst_ack_0,
          reqR => binary_2000_inst_req_1,
          ackR => binary_2000_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_2014_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_2009;
      tmp75_2015 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2014_inst_req_0,
          ackL => binary_2014_inst_ack_0,
          reqR => binary_2014_inst_req_1,
          ackR => binary_2014_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_2019_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp45_1931 & tmp40_1917;
      mask51_2020 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2019_inst_req_0,
          ackL => binary_2019_inst_ack_0,
          reqR => binary_2019_inst_req_1,
          ackR => binary_2019_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_2024_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask51_2020 & tmp50_1945;
      mask56_2025 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2024_inst_req_0,
          ackL => binary_2024_inst_ack_0,
          reqR => binary_2024_inst_req_1,
          ackR => binary_2024_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_2029_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask56_2025 & tmp55_1959;
      mask61x_xmaskedx_xmasked_2030 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2029_inst_req_0,
          ackL => binary_2029_inst_ack_0,
          reqR => binary_2029_inst_req_1,
          ackR => binary_2029_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_2034_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask61x_xmaskedx_xmasked_2030 & tmp60_1973;
      mask66x_xmaskedx_xmasked_2035 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2034_inst_req_0,
          ackL => binary_2034_inst_ack_0,
          reqR => binary_2034_inst_req_1,
          ackR => binary_2034_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_2039_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask66x_xmaskedx_xmasked_2035 & tmp65_1987;
      mask71x_xmasked_2040 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2039_inst_req_0,
          ackL => binary_2039_inst_ack_0,
          reqR => binary_2039_inst_req_1,
          ackR => binary_2039_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_2044_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask71x_xmasked_2040 & tmp70_2001;
      mask76_2045 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2044_inst_req_0,
          ackL => binary_2044_inst_ack_0,
          reqR => binary_2044_inst_req_1,
          ackR => binary_2044_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_2049_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask76_2045 & tmp75_2015;
      ins77_2050 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2049_inst_req_0,
          ackL => binary_2049_inst_ack_0,
          reqR => binary_2049_inst_req_1,
          ackR => binary_2049_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_2055_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_1816;
      exitcond_2056 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000011110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2055_inst_req_0,
          ackL => binary_2055_inst_ack_0,
          reqR => binary_2055_inst_req_1,
          ackR => binary_2055_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : binary_2087_inst 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_1816;
      indvarx_xnext_2088 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2087_inst_req_0,
          ackL => binary_2087_inst_ack_0,
          reqR => binary_2087_inst_req_1,
          ackR => binary_2087_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared load operator group (0) : ptr_deref_1626_load_0 ptr_deref_1912_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1626_load_0_req_0;
      reqL(0) <= ptr_deref_1912_load_0_req_0;
      ptr_deref_1626_load_0_ack_0 <= ackL(1);
      ptr_deref_1912_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1626_load_0_req_1;
      reqR(0) <= ptr_deref_1912_load_0_req_1;
      ptr_deref_1626_load_0_ack_1 <= ackR(1);
      ptr_deref_1912_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1626_word_address_0 & ptr_deref_1912_word_address_0;
      ptr_deref_1626_data_0 <= data_out(15 downto 8);
      ptr_deref_1912_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(7),
          mack => memory_space_0_lr_ack(7),
          maddr => memory_space_0_lr_addr(87 downto 77),
          mtag => memory_space_0_lr_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(7),
          mack => memory_space_0_lc_ack(7),
          mdata => memory_space_0_lc_data(63 downto 56),
          mtag => memory_space_0_lc_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1920_load_0 ptr_deref_1639_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1920_load_0_req_0;
      reqL(0) <= ptr_deref_1639_load_0_req_0;
      ptr_deref_1920_load_0_ack_0 <= ackL(1);
      ptr_deref_1639_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1920_load_0_req_1;
      reqR(0) <= ptr_deref_1639_load_0_req_1;
      ptr_deref_1920_load_0_ack_1 <= ackR(1);
      ptr_deref_1639_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1920_word_address_0 & ptr_deref_1639_word_address_0;
      ptr_deref_1920_data_0 <= data_out(15 downto 8);
      ptr_deref_1639_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(6),
          mack => memory_space_0_lr_ack(6),
          maddr => memory_space_0_lr_addr(76 downto 66),
          mtag => memory_space_0_lr_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(6),
          mack => memory_space_0_lc_ack(6),
          mdata => memory_space_0_lc_data(55 downto 48),
          mtag => memory_space_0_lc_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1934_load_0 ptr_deref_1658_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1934_load_0_req_0;
      reqL(0) <= ptr_deref_1658_load_0_req_0;
      ptr_deref_1934_load_0_ack_0 <= ackL(1);
      ptr_deref_1658_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1934_load_0_req_1;
      reqR(0) <= ptr_deref_1658_load_0_req_1;
      ptr_deref_1934_load_0_ack_1 <= ackR(1);
      ptr_deref_1658_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1934_word_address_0 & ptr_deref_1658_word_address_0;
      ptr_deref_1934_data_0 <= data_out(15 downto 8);
      ptr_deref_1658_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(5),
          mack => memory_space_0_lr_ack(5),
          maddr => memory_space_0_lr_addr(65 downto 55),
          mtag => memory_space_0_lr_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(5),
          mack => memory_space_0_lc_ack(5),
          mdata => memory_space_0_lc_data(47 downto 40),
          mtag => memory_space_0_lc_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1677_load_0 ptr_deref_1948_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1677_load_0_req_0;
      reqL(0) <= ptr_deref_1948_load_0_req_0;
      ptr_deref_1677_load_0_ack_0 <= ackL(1);
      ptr_deref_1948_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1677_load_0_req_1;
      reqR(0) <= ptr_deref_1948_load_0_req_1;
      ptr_deref_1677_load_0_ack_1 <= ackR(1);
      ptr_deref_1948_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1677_word_address_0 & ptr_deref_1948_word_address_0;
      ptr_deref_1677_data_0 <= data_out(15 downto 8);
      ptr_deref_1948_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(4),
          mack => memory_space_0_lr_ack(4),
          maddr => memory_space_0_lr_addr(54 downto 44),
          mtag => memory_space_0_lr_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(4),
          mack => memory_space_0_lc_ack(4),
          mdata => memory_space_0_lc_data(39 downto 32),
          mtag => memory_space_0_lc_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1696_load_0 ptr_deref_1962_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1696_load_0_req_0;
      reqL(0) <= ptr_deref_1962_load_0_req_0;
      ptr_deref_1696_load_0_ack_0 <= ackL(1);
      ptr_deref_1962_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1696_load_0_req_1;
      reqR(0) <= ptr_deref_1962_load_0_req_1;
      ptr_deref_1696_load_0_ack_1 <= ackR(1);
      ptr_deref_1962_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1696_word_address_0 & ptr_deref_1962_word_address_0;
      ptr_deref_1696_data_0 <= data_out(15 downto 8);
      ptr_deref_1962_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(3),
          mack => memory_space_0_lr_ack(3),
          maddr => memory_space_0_lr_addr(43 downto 33),
          mtag => memory_space_0_lr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(3),
          mack => memory_space_0_lc_ack(3),
          mdata => memory_space_0_lc_data(31 downto 24),
          mtag => memory_space_0_lc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1715_load_0 ptr_deref_1976_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1715_load_0_req_0;
      reqL(0) <= ptr_deref_1976_load_0_req_0;
      ptr_deref_1715_load_0_ack_0 <= ackL(1);
      ptr_deref_1976_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1715_load_0_req_1;
      reqR(0) <= ptr_deref_1976_load_0_req_1;
      ptr_deref_1715_load_0_ack_1 <= ackR(1);
      ptr_deref_1976_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1715_word_address_0 & ptr_deref_1976_word_address_0;
      ptr_deref_1715_data_0 <= data_out(15 downto 8);
      ptr_deref_1976_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(2),
          mack => memory_space_0_lr_ack(2),
          maddr => memory_space_0_lr_addr(32 downto 22),
          mtag => memory_space_0_lr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(2),
          mack => memory_space_0_lc_ack(2),
          mdata => memory_space_0_lc_data(23 downto 16),
          mtag => memory_space_0_lc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_1729_load_0 ptr_deref_1990_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1729_load_0_req_0;
      reqL(0) <= ptr_deref_1990_load_0_req_0;
      ptr_deref_1729_load_0_ack_0 <= ackL(1);
      ptr_deref_1990_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1729_load_0_req_1;
      reqR(0) <= ptr_deref_1990_load_0_req_1;
      ptr_deref_1729_load_0_ack_1 <= ackR(1);
      ptr_deref_1990_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1729_word_address_0 & ptr_deref_1990_word_address_0;
      ptr_deref_1729_data_0 <= data_out(15 downto 8);
      ptr_deref_1990_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(1),
          mack => memory_space_0_lr_ack(1),
          maddr => memory_space_0_lr_addr(21 downto 11),
          mtag => memory_space_0_lr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(1),
          mack => memory_space_0_lc_ack(1),
          mdata => memory_space_0_lc_data(15 downto 8),
          mtag => memory_space_0_lc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_1748_load_0 ptr_deref_2004_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1748_load_0_req_0;
      reqL(0) <= ptr_deref_2004_load_0_req_0;
      ptr_deref_1748_load_0_ack_0 <= ackL(1);
      ptr_deref_2004_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1748_load_0_req_1;
      reqR(0) <= ptr_deref_2004_load_0_req_1;
      ptr_deref_1748_load_0_ack_1 <= ackR(1);
      ptr_deref_2004_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1748_word_address_0 & ptr_deref_2004_word_address_0;
      ptr_deref_1748_data_0 <= data_out(15 downto 8);
      ptr_deref_2004_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(10 downto 0),
          mtag => memory_space_0_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(7 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared inport operator group (0) : simple_obj_ref_1613_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1613_inst_req_0;
      simple_obj_ref_1613_inst_ack_0 <= ack(0);
      tmp_1614 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => midpipe_pipe_read_req(0),
          oack => midpipe_pipe_read_ack(0),
          odata => midpipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : simple_obj_ref_1801_inst simple_obj_ref_2091_inst simple_obj_ref_2070_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_1801_inst_req_0;
      req(1) <= simple_obj_ref_2091_inst_req_0;
      req(0) <= simple_obj_ref_2070_inst_req_0;
      simple_obj_ref_1801_inst_ack_0 <= ack(2);
      simple_obj_ref_2091_inst_ack_0 <= ack(1);
      simple_obj_ref_2070_inst_ack_0 <= ack(0);
      data_in <= type_cast_1803_wire_constant & type_cast_2093_wire_constant & type_cast_2072_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 3,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_ctrl_pipe_write_req(0),
          oack => out_ctrl_pipe_write_ack(0),
          odata => out_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_1811_inst simple_obj_ref_2101_inst simple_obj_ref_2080_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_1811_inst_req_0;
      req(1) <= simple_obj_ref_2101_inst_req_0;
      req(0) <= simple_obj_ref_2080_inst_req_0;
      simple_obj_ref_1811_inst_ack_0 <= ack(2);
      simple_obj_ref_2101_inst_ack_0 <= ack(1);
      simple_obj_ref_2080_inst_ack_0 <= ack(0);
      data_in <= ins38_1794 & ins77_2050 & ins77_2050;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 3,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_2110_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2110_inst_req_0;
      simple_obj_ref_2110_inst_ack_0 <= ack(0);
      data_in <= type_cast_2112_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : simple_obj_ref_2120_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2120_inst_req_0;
      simple_obj_ref_2120_inst_ack_0 <= ack(0);
      data_in <= tmp_1614;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_put_pipe_write_req(0),
          oack => free_queue_put_pipe_write_ack(0),
          odata => free_queue_put_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_ctrl_pipe_write_data: in std_logic_vector(7 downto 0);
    in_ctrl_pipe_write_req : in std_logic_vector(0 downto 0);
    in_ctrl_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_pipe_write_data: in std_logic_vector(63 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_data: out std_logic_vector(7 downto 0);
    out_ctrl_pipe_read_req : in std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(63 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(7 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(7 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(87 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(15 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(7 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(7 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(15 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(8 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(8 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(98 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(71 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(8 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(8 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(17 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(7 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_10
  signal memory_space_10_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_10_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_10_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_10_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_11
  signal memory_space_11_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_11_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_11_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_11_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(14 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(39 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(9 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(9 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_9
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module default_initializer_foo
  component default_initializer_foo is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_foo
  signal default_initializer_foo_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_foo_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_foo_start_req : std_logic;
  signal default_initializer_foo_start_ack : std_logic;
  signal default_initializer_foo_fin_req   : std_logic;
  signal default_initializer_foo_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_foo
  signal default_initializer_foo_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_foo_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_foo_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_foo_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_foo_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_foo_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_free_queue
  component default_initializer_free_queue is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_free_queue
  signal default_initializer_free_queue_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_free_queue_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_start_req : std_logic;
  signal default_initializer_free_queue_start_ack : std_logic;
  signal default_initializer_free_queue_fin_req   : std_logic;
  signal default_initializer_free_queue_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_free_queue
  signal default_initializer_free_queue_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_free_queue_ram
  component default_initializer_free_queue_ram is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_free_queue_ram
  signal default_initializer_free_queue_ram_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_free_queue_ram_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_start_req : std_logic;
  signal default_initializer_free_queue_ram_start_ack : std_logic;
  signal default_initializer_free_queue_ram_fin_req   : std_logic;
  signal default_initializer_free_queue_ram_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_free_queue_ram
  signal default_initializer_free_queue_ram_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_free_queue_ram_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr
  component default_initializer_xx_xstr is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(4 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr
  signal default_initializer_xx_xstr_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_start_req : std_logic;
  signal default_initializer_xx_xstr_start_ack : std_logic;
  signal default_initializer_xx_xstr_fin_req   : std_logic;
  signal default_initializer_xx_xstr_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr
  signal default_initializer_xx_xstr_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr1
  component default_initializer_xx_xstr1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr1
  signal default_initializer_xx_xstr1_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr1_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_start_req : std_logic;
  signal default_initializer_xx_xstr1_start_ack : std_logic;
  signal default_initializer_xx_xstr1_fin_req   : std_logic;
  signal default_initializer_xx_xstr1_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr1
  signal default_initializer_xx_xstr1_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr1_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr2
  component default_initializer_xx_xstr2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr2
  signal default_initializer_xx_xstr2_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr2_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_start_req : std_logic;
  signal default_initializer_xx_xstr2_start_ack : std_logic;
  signal default_initializer_xx_xstr2_fin_req   : std_logic;
  signal default_initializer_xx_xstr2_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr2
  signal default_initializer_xx_xstr2_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr2_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr3
  component default_initializer_xx_xstr3 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr3
  signal default_initializer_xx_xstr3_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr3_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_start_req : std_logic;
  signal default_initializer_xx_xstr3_start_ack : std_logic;
  signal default_initializer_xx_xstr3_fin_req   : std_logic;
  signal default_initializer_xx_xstr3_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr3
  signal default_initializer_xx_xstr3_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr3_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr4
  component default_initializer_xx_xstr4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr4
  signal default_initializer_xx_xstr4_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr4_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_start_req : std_logic;
  signal default_initializer_xx_xstr4_start_ack : std_logic;
  signal default_initializer_xx_xstr4_fin_req   : std_logic;
  signal default_initializer_xx_xstr4_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr4
  signal default_initializer_xx_xstr4_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr5
  component default_initializer_xx_xstr5 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr5
  signal default_initializer_xx_xstr5_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr5_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_start_req : std_logic;
  signal default_initializer_xx_xstr5_start_ack : std_logic;
  signal default_initializer_xx_xstr5_fin_req   : std_logic;
  signal default_initializer_xx_xstr5_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr5
  signal default_initializer_xx_xstr5_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr5_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr6
  component default_initializer_xx_xstr6 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_9_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_9_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_9_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_9_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_9_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_9_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr6
  signal default_initializer_xx_xstr6_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr6_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_start_req : std_logic;
  signal default_initializer_xx_xstr6_start_ack : std_logic;
  signal default_initializer_xx_xstr6_fin_req   : std_logic;
  signal default_initializer_xx_xstr6_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr6
  signal default_initializer_xx_xstr6_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr6_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr7
  component default_initializer_xx_xstr7 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_10_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_10_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_10_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_10_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_10_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_10_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr7
  signal default_initializer_xx_xstr7_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr7_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_start_req : std_logic;
  signal default_initializer_xx_xstr7_start_ack : std_logic;
  signal default_initializer_xx_xstr7_fin_req   : std_logic;
  signal default_initializer_xx_xstr7_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr7
  signal default_initializer_xx_xstr7_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr7_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module default_initializer_xx_xstr8
  component default_initializer_xx_xstr8 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_11_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_11_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_11_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_11_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_11_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_11_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module default_initializer_xx_xstr8
  signal default_initializer_xx_xstr8_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal default_initializer_xx_xstr8_tag_out   : std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_start_req : std_logic;
  signal default_initializer_xx_xstr8_start_ack : std_logic;
  signal default_initializer_xx_xstr8_fin_req   : std_logic;
  signal default_initializer_xx_xstr8_fin_ack : std_logic;
  -- caller side aggregated signals for module default_initializer_xx_xstr8
  signal default_initializer_xx_xstr8_call_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_call_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_return_reqs: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_return_acks: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_call_tag: std_logic_vector(0 downto 0);
  signal default_initializer_xx_xstr8_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module free_queue_manager
  component free_queue_manager is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(3 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(3 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(3 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(3 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(7 downto 0);
      free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_ack_pipe_write_data : out  std_logic_vector(7 downto 0);
      free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
      global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module free_queue_manager
  signal free_queue_manager_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal free_queue_manager_tag_out   : std_logic_vector(0 downto 0);
  signal free_queue_manager_start_req : std_logic;
  signal free_queue_manager_start_ack : std_logic;
  signal free_queue_manager_fin_req   : std_logic;
  signal free_queue_manager_fin_ack : std_logic;
  -- declarations related to module global_storage_initializer_x
  component global_storage_initializer_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      default_initializer_xx_xstr2_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr2_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr4_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_foo_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_foo_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_foo_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_foo_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_foo_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_foo_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_free_queue_ram_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr5_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr8_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr7_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr1_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr3_return_tag :  in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_call_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_call_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_call_tag  :  out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_return_reqs : out  std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_return_acks : in   std_logic_vector(0 downto 0);
      default_initializer_xx_xstr6_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module global_storage_initializer_x
  signal global_storage_initializer_x_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal global_storage_initializer_x_tag_out   : std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_start_req : std_logic;
  signal global_storage_initializer_x_start_ack : std_logic;
  signal global_storage_initializer_x_fin_req   : std_logic;
  signal global_storage_initializer_x_fin_ack : std_logic;
  -- caller side aggregated signals for module global_storage_initializer_x
  signal global_storage_initializer_x_call_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_tag: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module wrapper_input
  component wrapper_input is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_0_sr_req : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(7 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(87 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(15 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(7 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(7 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(15 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
      in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      midpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      midpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      midpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_input
  signal wrapper_input_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_input_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_input_start_req : std_logic;
  signal wrapper_input_start_ack : std_logic;
  signal wrapper_input_fin_req   : std_logic;
  signal wrapper_input_fin_ack : std_logic;
  -- declarations related to module wrapper_output
  component wrapper_output is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_0_lr_req : out  std_logic_vector(7 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(7 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(87 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(15 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(7 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(7 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(15 downto 0);
      midpipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      midpipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      midpipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
      out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_output
  signal wrapper_output_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_output_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_output_start_req : std_logic;
  signal wrapper_output_start_ack : std_logic;
  signal wrapper_output_fin_req   : std_logic;
  signal wrapper_output_fin_ack : std_logic;
  -- aggregate signals for write to pipe free_queue_ack
  signal free_queue_ack_pipe_write_data: std_logic_vector(7 downto 0);
  signal free_queue_ack_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_ack_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_ack
  signal free_queue_ack_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_ack_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_ack_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_get
  signal free_queue_get_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_get
  signal free_queue_get_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_put
  signal free_queue_put_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_put
  signal free_queue_put_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_request
  signal free_queue_request_pipe_write_data: std_logic_vector(15 downto 0);
  signal free_queue_request_pipe_write_req: std_logic_vector(1 downto 0);
  signal free_queue_request_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe free_queue_request
  signal free_queue_request_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_request_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_request_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_ctrl
  signal in_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal in_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe midpipe
  signal midpipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal midpipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal midpipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe midpipe
  signal midpipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal midpipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal midpipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_ctrl
  signal out_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal out_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module default_initializer_foo
  -- call arbiter for module default_initializer_foo
  default_initializer_foo_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_foo_call_reqs,
      call_acks => default_initializer_foo_call_acks,
      return_reqs => default_initializer_foo_return_reqs,
      return_acks => default_initializer_foo_return_acks,
      call_tag  => default_initializer_foo_call_tag,
      return_tag  => default_initializer_foo_return_tag,
      call_mtag => default_initializer_foo_tag_in,
      return_mtag => default_initializer_foo_tag_out,
      call_mreq => default_initializer_foo_start_req,
      call_mack => default_initializer_foo_start_ack,
      return_mreq => default_initializer_foo_fin_req,
      return_mack => default_initializer_foo_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_foo_instance:default_initializer_foo-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_foo_start_req,
      start_ack => default_initializer_foo_start_ack,
      fin_req => default_initializer_foo_fin_req,
      fin_ack => default_initializer_foo_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(1 downto 1),
      memory_space_1_sr_ack => memory_space_1_sr_ack(1 downto 1),
      memory_space_1_sr_addr => memory_space_1_sr_addr(7 downto 4),
      memory_space_1_sr_data => memory_space_1_sr_data(15 downto 8),
      memory_space_1_sr_tag => memory_space_1_sr_tag(1 downto 1),
      memory_space_1_sc_req => memory_space_1_sc_req(1 downto 1),
      memory_space_1_sc_ack => memory_space_1_sc_ack(1 downto 1),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 1),
      tag_in => default_initializer_foo_tag_in,
      tag_out => default_initializer_foo_tag_out-- 
    ); -- 
  -- module default_initializer_free_queue
  -- call arbiter for module default_initializer_free_queue
  default_initializer_free_queue_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_free_queue_call_reqs,
      call_acks => default_initializer_free_queue_call_acks,
      return_reqs => default_initializer_free_queue_return_reqs,
      return_acks => default_initializer_free_queue_return_acks,
      call_tag  => default_initializer_free_queue_call_tag,
      return_tag  => default_initializer_free_queue_return_tag,
      call_mtag => default_initializer_free_queue_tag_in,
      return_mtag => default_initializer_free_queue_tag_out,
      call_mreq => default_initializer_free_queue_start_req,
      call_mack => default_initializer_free_queue_start_ack,
      return_mreq => default_initializer_free_queue_fin_req,
      return_mack => default_initializer_free_queue_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_free_queue_instance:default_initializer_free_queue-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_free_queue_start_req,
      start_ack => default_initializer_free_queue_start_ack,
      fin_req => default_initializer_free_queue_fin_req,
      fin_ack => default_initializer_free_queue_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(4 downto 4),
      memory_space_2_sr_ack => memory_space_2_sr_ack(4 downto 4),
      memory_space_2_sr_addr => memory_space_2_sr_addr(14 downto 12),
      memory_space_2_sr_data => memory_space_2_sr_data(39 downto 32),
      memory_space_2_sr_tag => memory_space_2_sr_tag(9 downto 8),
      memory_space_2_sc_req => memory_space_2_sc_req(4 downto 4),
      memory_space_2_sc_ack => memory_space_2_sc_ack(4 downto 4),
      memory_space_2_sc_tag => memory_space_2_sc_tag(9 downto 8),
      tag_in => default_initializer_free_queue_tag_in,
      tag_out => default_initializer_free_queue_tag_out-- 
    ); -- 
  -- module default_initializer_free_queue_ram
  -- call arbiter for module default_initializer_free_queue_ram
  default_initializer_free_queue_ram_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_free_queue_ram_call_reqs,
      call_acks => default_initializer_free_queue_ram_call_acks,
      return_reqs => default_initializer_free_queue_ram_return_reqs,
      return_acks => default_initializer_free_queue_ram_return_acks,
      call_tag  => default_initializer_free_queue_ram_call_tag,
      return_tag  => default_initializer_free_queue_ram_return_tag,
      call_mtag => default_initializer_free_queue_ram_tag_in,
      return_mtag => default_initializer_free_queue_ram_tag_out,
      call_mreq => default_initializer_free_queue_ram_start_req,
      call_mack => default_initializer_free_queue_ram_start_ack,
      return_mreq => default_initializer_free_queue_ram_fin_req,
      return_mack => default_initializer_free_queue_ram_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_free_queue_ram_instance:default_initializer_free_queue_ram-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_free_queue_ram_start_req,
      start_ack => default_initializer_free_queue_ram_start_ack,
      fin_req => default_initializer_free_queue_ram_fin_req,
      fin_ack => default_initializer_free_queue_ram_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(8 downto 8),
      memory_space_0_sr_ack => memory_space_0_sr_ack(8 downto 8),
      memory_space_0_sr_addr => memory_space_0_sr_addr(98 downto 88),
      memory_space_0_sr_data => memory_space_0_sr_data(71 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 16),
      memory_space_0_sc_req => memory_space_0_sc_req(8 downto 8),
      memory_space_0_sc_ack => memory_space_0_sc_ack(8 downto 8),
      memory_space_0_sc_tag => memory_space_0_sc_tag(17 downto 16),
      tag_in => default_initializer_free_queue_ram_tag_in,
      tag_out => default_initializer_free_queue_ram_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr
  -- call arbiter for module default_initializer_xx_xstr
  default_initializer_xx_xstr_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr_call_reqs,
      call_acks => default_initializer_xx_xstr_call_acks,
      return_reqs => default_initializer_xx_xstr_return_reqs,
      return_acks => default_initializer_xx_xstr_return_acks,
      call_tag  => default_initializer_xx_xstr_call_tag,
      return_tag  => default_initializer_xx_xstr_return_tag,
      call_mtag => default_initializer_xx_xstr_tag_in,
      return_mtag => default_initializer_xx_xstr_tag_out,
      call_mreq => default_initializer_xx_xstr_start_req,
      call_mack => default_initializer_xx_xstr_start_ack,
      return_mreq => default_initializer_xx_xstr_fin_req,
      return_mack => default_initializer_xx_xstr_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr_instance:default_initializer_xx_xstr-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr_start_req,
      start_ack => default_initializer_xx_xstr_start_ack,
      fin_req => default_initializer_xx_xstr_fin_req,
      fin_ack => default_initializer_xx_xstr_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(4 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(7 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(4 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 0),
      tag_in => default_initializer_xx_xstr_tag_in,
      tag_out => default_initializer_xx_xstr_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr1
  -- call arbiter for module default_initializer_xx_xstr1
  default_initializer_xx_xstr1_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr1_call_reqs,
      call_acks => default_initializer_xx_xstr1_call_acks,
      return_reqs => default_initializer_xx_xstr1_return_reqs,
      return_acks => default_initializer_xx_xstr1_return_acks,
      call_tag  => default_initializer_xx_xstr1_call_tag,
      return_tag  => default_initializer_xx_xstr1_return_tag,
      call_mtag => default_initializer_xx_xstr1_tag_in,
      return_mtag => default_initializer_xx_xstr1_tag_out,
      call_mreq => default_initializer_xx_xstr1_start_req,
      call_mack => default_initializer_xx_xstr1_start_ack,
      return_mreq => default_initializer_xx_xstr1_fin_req,
      return_mack => default_initializer_xx_xstr1_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr1_instance:default_initializer_xx_xstr1-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr1_start_req,
      start_ack => default_initializer_xx_xstr1_start_ack,
      fin_req => default_initializer_xx_xstr1_fin_req,
      fin_ack => default_initializer_xx_xstr1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(3 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(7 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(3 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr1_tag_in,
      tag_out => default_initializer_xx_xstr1_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr2
  -- call arbiter for module default_initializer_xx_xstr2
  default_initializer_xx_xstr2_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr2_call_reqs,
      call_acks => default_initializer_xx_xstr2_call_acks,
      return_reqs => default_initializer_xx_xstr2_return_reqs,
      return_acks => default_initializer_xx_xstr2_return_acks,
      call_tag  => default_initializer_xx_xstr2_call_tag,
      return_tag  => default_initializer_xx_xstr2_return_tag,
      call_mtag => default_initializer_xx_xstr2_tag_in,
      return_mtag => default_initializer_xx_xstr2_tag_out,
      call_mreq => default_initializer_xx_xstr2_start_req,
      call_mack => default_initializer_xx_xstr2_start_ack,
      return_mreq => default_initializer_xx_xstr2_fin_req,
      return_mack => default_initializer_xx_xstr2_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr2_instance:default_initializer_xx_xstr2-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr2_start_req,
      start_ack => default_initializer_xx_xstr2_start_ack,
      fin_req => default_initializer_xx_xstr2_fin_req,
      fin_ack => default_initializer_xx_xstr2_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(3 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(7 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(3 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr2_tag_in,
      tag_out => default_initializer_xx_xstr2_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr3
  -- call arbiter for module default_initializer_xx_xstr3
  default_initializer_xx_xstr3_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr3_call_reqs,
      call_acks => default_initializer_xx_xstr3_call_acks,
      return_reqs => default_initializer_xx_xstr3_return_reqs,
      return_acks => default_initializer_xx_xstr3_return_acks,
      call_tag  => default_initializer_xx_xstr3_call_tag,
      return_tag  => default_initializer_xx_xstr3_return_tag,
      call_mtag => default_initializer_xx_xstr3_tag_in,
      return_mtag => default_initializer_xx_xstr3_tag_out,
      call_mreq => default_initializer_xx_xstr3_start_req,
      call_mack => default_initializer_xx_xstr3_start_ack,
      return_mreq => default_initializer_xx_xstr3_fin_req,
      return_mack => default_initializer_xx_xstr3_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr3_instance:default_initializer_xx_xstr3-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr3_start_req,
      start_ack => default_initializer_xx_xstr3_start_ack,
      fin_req => default_initializer_xx_xstr3_fin_req,
      fin_ack => default_initializer_xx_xstr3_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(3 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(7 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(3 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr3_tag_in,
      tag_out => default_initializer_xx_xstr3_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr4
  -- call arbiter for module default_initializer_xx_xstr4
  default_initializer_xx_xstr4_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr4_call_reqs,
      call_acks => default_initializer_xx_xstr4_call_acks,
      return_reqs => default_initializer_xx_xstr4_return_reqs,
      return_acks => default_initializer_xx_xstr4_return_acks,
      call_tag  => default_initializer_xx_xstr4_call_tag,
      return_tag  => default_initializer_xx_xstr4_return_tag,
      call_mtag => default_initializer_xx_xstr4_tag_in,
      return_mtag => default_initializer_xx_xstr4_tag_out,
      call_mreq => default_initializer_xx_xstr4_start_req,
      call_mack => default_initializer_xx_xstr4_start_ack,
      return_mreq => default_initializer_xx_xstr4_fin_req,
      return_mack => default_initializer_xx_xstr4_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr4_instance:default_initializer_xx_xstr4-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr4_start_req,
      start_ack => default_initializer_xx_xstr4_start_ack,
      fin_req => default_initializer_xx_xstr4_fin_req,
      fin_ack => default_initializer_xx_xstr4_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(3 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(7 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(3 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr4_tag_in,
      tag_out => default_initializer_xx_xstr4_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr5
  -- call arbiter for module default_initializer_xx_xstr5
  default_initializer_xx_xstr5_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr5_call_reqs,
      call_acks => default_initializer_xx_xstr5_call_acks,
      return_reqs => default_initializer_xx_xstr5_return_reqs,
      return_acks => default_initializer_xx_xstr5_return_acks,
      call_tag  => default_initializer_xx_xstr5_call_tag,
      return_tag  => default_initializer_xx_xstr5_return_tag,
      call_mtag => default_initializer_xx_xstr5_tag_in,
      return_mtag => default_initializer_xx_xstr5_tag_out,
      call_mreq => default_initializer_xx_xstr5_start_req,
      call_mack => default_initializer_xx_xstr5_start_ack,
      return_mreq => default_initializer_xx_xstr5_fin_req,
      return_mack => default_initializer_xx_xstr5_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr5_instance:default_initializer_xx_xstr5-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr5_start_req,
      start_ack => default_initializer_xx_xstr5_start_ack,
      fin_req => default_initializer_xx_xstr5_fin_req,
      fin_ack => default_initializer_xx_xstr5_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(3 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(7 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(3 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr5_tag_in,
      tag_out => default_initializer_xx_xstr5_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr6
  -- call arbiter for module default_initializer_xx_xstr6
  default_initializer_xx_xstr6_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr6_call_reqs,
      call_acks => default_initializer_xx_xstr6_call_acks,
      return_reqs => default_initializer_xx_xstr6_return_reqs,
      return_acks => default_initializer_xx_xstr6_return_acks,
      call_tag  => default_initializer_xx_xstr6_call_tag,
      return_tag  => default_initializer_xx_xstr6_return_tag,
      call_mtag => default_initializer_xx_xstr6_tag_in,
      return_mtag => default_initializer_xx_xstr6_tag_out,
      call_mreq => default_initializer_xx_xstr6_start_req,
      call_mack => default_initializer_xx_xstr6_start_ack,
      return_mreq => default_initializer_xx_xstr6_fin_req,
      return_mack => default_initializer_xx_xstr6_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr6_instance:default_initializer_xx_xstr6-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr6_start_req,
      start_ack => default_initializer_xx_xstr6_start_ack,
      fin_req => default_initializer_xx_xstr6_fin_req,
      fin_ack => default_initializer_xx_xstr6_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_9_sr_req => memory_space_9_sr_req(0 downto 0),
      memory_space_9_sr_ack => memory_space_9_sr_ack(0 downto 0),
      memory_space_9_sr_addr => memory_space_9_sr_addr(3 downto 0),
      memory_space_9_sr_data => memory_space_9_sr_data(7 downto 0),
      memory_space_9_sr_tag => memory_space_9_sr_tag(3 downto 0),
      memory_space_9_sc_req => memory_space_9_sc_req(0 downto 0),
      memory_space_9_sc_ack => memory_space_9_sc_ack(0 downto 0),
      memory_space_9_sc_tag => memory_space_9_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr6_tag_in,
      tag_out => default_initializer_xx_xstr6_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr7
  -- call arbiter for module default_initializer_xx_xstr7
  default_initializer_xx_xstr7_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr7_call_reqs,
      call_acks => default_initializer_xx_xstr7_call_acks,
      return_reqs => default_initializer_xx_xstr7_return_reqs,
      return_acks => default_initializer_xx_xstr7_return_acks,
      call_tag  => default_initializer_xx_xstr7_call_tag,
      return_tag  => default_initializer_xx_xstr7_return_tag,
      call_mtag => default_initializer_xx_xstr7_tag_in,
      return_mtag => default_initializer_xx_xstr7_tag_out,
      call_mreq => default_initializer_xx_xstr7_start_req,
      call_mack => default_initializer_xx_xstr7_start_ack,
      return_mreq => default_initializer_xx_xstr7_fin_req,
      return_mack => default_initializer_xx_xstr7_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr7_instance:default_initializer_xx_xstr7-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr7_start_req,
      start_ack => default_initializer_xx_xstr7_start_ack,
      fin_req => default_initializer_xx_xstr7_fin_req,
      fin_ack => default_initializer_xx_xstr7_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_10_sr_req => memory_space_10_sr_req(0 downto 0),
      memory_space_10_sr_ack => memory_space_10_sr_ack(0 downto 0),
      memory_space_10_sr_addr => memory_space_10_sr_addr(3 downto 0),
      memory_space_10_sr_data => memory_space_10_sr_data(7 downto 0),
      memory_space_10_sr_tag => memory_space_10_sr_tag(3 downto 0),
      memory_space_10_sc_req => memory_space_10_sc_req(0 downto 0),
      memory_space_10_sc_ack => memory_space_10_sc_ack(0 downto 0),
      memory_space_10_sc_tag => memory_space_10_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr7_tag_in,
      tag_out => default_initializer_xx_xstr7_tag_out-- 
    ); -- 
  -- module default_initializer_xx_xstr8
  -- call arbiter for module default_initializer_xx_xstr8
  default_initializer_xx_xstr8_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => default_initializer_xx_xstr8_call_reqs,
      call_acks => default_initializer_xx_xstr8_call_acks,
      return_reqs => default_initializer_xx_xstr8_return_reqs,
      return_acks => default_initializer_xx_xstr8_return_acks,
      call_tag  => default_initializer_xx_xstr8_call_tag,
      return_tag  => default_initializer_xx_xstr8_return_tag,
      call_mtag => default_initializer_xx_xstr8_tag_in,
      return_mtag => default_initializer_xx_xstr8_tag_out,
      call_mreq => default_initializer_xx_xstr8_start_req,
      call_mack => default_initializer_xx_xstr8_start_ack,
      return_mreq => default_initializer_xx_xstr8_fin_req,
      return_mack => default_initializer_xx_xstr8_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  default_initializer_xx_xstr8_instance:default_initializer_xx_xstr8-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => default_initializer_xx_xstr8_start_req,
      start_ack => default_initializer_xx_xstr8_start_ack,
      fin_req => default_initializer_xx_xstr8_fin_req,
      fin_ack => default_initializer_xx_xstr8_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_11_sr_req => memory_space_11_sr_req(0 downto 0),
      memory_space_11_sr_ack => memory_space_11_sr_ack(0 downto 0),
      memory_space_11_sr_addr => memory_space_11_sr_addr(3 downto 0),
      memory_space_11_sr_data => memory_space_11_sr_data(7 downto 0),
      memory_space_11_sr_tag => memory_space_11_sr_tag(3 downto 0),
      memory_space_11_sc_req => memory_space_11_sc_req(0 downto 0),
      memory_space_11_sc_ack => memory_space_11_sc_ack(0 downto 0),
      memory_space_11_sc_tag => memory_space_11_sc_tag(3 downto 0),
      tag_in => default_initializer_xx_xstr8_tag_in,
      tag_out => default_initializer_xx_xstr8_tag_out-- 
    ); -- 
  -- module free_queue_manager
  free_queue_manager_instance:free_queue_manager-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => free_queue_manager_start_req,
      start_ack => free_queue_manager_start_ack,
      fin_req => free_queue_manager_fin_req,
      fin_ack => free_queue_manager_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(2 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(1 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(7 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(11 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(7 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(7 downto 0),
      free_queue_request_pipe_read_req => free_queue_request_pipe_read_req(0 downto 0),
      free_queue_request_pipe_read_ack => free_queue_request_pipe_read_ack(0 downto 0),
      free_queue_request_pipe_read_data => free_queue_request_pipe_read_data(7 downto 0),
      free_queue_put_pipe_read_req => free_queue_put_pipe_read_req(0 downto 0),
      free_queue_put_pipe_read_ack => free_queue_put_pipe_read_ack(0 downto 0),
      free_queue_put_pipe_read_data => free_queue_put_pipe_read_data(31 downto 0),
      free_queue_ack_pipe_write_req => free_queue_ack_pipe_write_req(0 downto 0),
      free_queue_ack_pipe_write_ack => free_queue_ack_pipe_write_ack(0 downto 0),
      free_queue_ack_pipe_write_data => free_queue_ack_pipe_write_data(7 downto 0),
      free_queue_get_pipe_write_req => free_queue_get_pipe_write_req(0 downto 0),
      free_queue_get_pipe_write_ack => free_queue_get_pipe_write_ack(0 downto 0),
      free_queue_get_pipe_write_data => free_queue_get_pipe_write_data(31 downto 0),
      global_storage_initializer_x_call_reqs => global_storage_initializer_x_call_reqs(0 downto 0),
      global_storage_initializer_x_call_acks => global_storage_initializer_x_call_acks(0 downto 0),
      global_storage_initializer_x_call_tag => global_storage_initializer_x_call_tag(0 downto 0),
      global_storage_initializer_x_return_reqs => global_storage_initializer_x_return_reqs(0 downto 0),
      global_storage_initializer_x_return_acks => global_storage_initializer_x_return_acks(0 downto 0),
      global_storage_initializer_x_return_tag => global_storage_initializer_x_return_tag(0 downto 0),
      tag_in => free_queue_manager_tag_in,
      tag_out => free_queue_manager_tag_out-- 
    ); -- 
  -- module will be run forever 
  free_queue_manager_tag_in <= (others => '0');
  free_queue_manager_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => free_queue_manager_start_req, start_ack => free_queue_manager_start_ack,  fin_req => free_queue_manager_fin_req,  fin_ack => free_queue_manager_fin_ack);
  -- module global_storage_initializer_x
  -- call arbiter for module global_storage_initializer_x
  global_storage_initializer_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => global_storage_initializer_x_call_reqs,
      call_acks => global_storage_initializer_x_call_acks,
      return_reqs => global_storage_initializer_x_return_reqs,
      return_acks => global_storage_initializer_x_return_acks,
      call_tag  => global_storage_initializer_x_call_tag,
      return_tag  => global_storage_initializer_x_return_tag,
      call_mtag => global_storage_initializer_x_tag_in,
      return_mtag => global_storage_initializer_x_tag_out,
      call_mreq => global_storage_initializer_x_start_req,
      call_mack => global_storage_initializer_x_start_ack,
      return_mreq => global_storage_initializer_x_fin_req,
      return_mack => global_storage_initializer_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  global_storage_initializer_x_instance:global_storage_initializer_x-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => global_storage_initializer_x_start_req,
      start_ack => global_storage_initializer_x_start_ack,
      fin_req => global_storage_initializer_x_fin_req,
      fin_ack => global_storage_initializer_x_fin_ack,
      clk => clk,
      reset => reset,
      default_initializer_foo_call_reqs => default_initializer_foo_call_reqs(0 downto 0),
      default_initializer_foo_call_acks => default_initializer_foo_call_acks(0 downto 0),
      default_initializer_foo_call_tag => default_initializer_foo_call_tag(0 downto 0),
      default_initializer_foo_return_reqs => default_initializer_foo_return_reqs(0 downto 0),
      default_initializer_foo_return_acks => default_initializer_foo_return_acks(0 downto 0),
      default_initializer_foo_return_tag => default_initializer_foo_return_tag(0 downto 0),
      default_initializer_free_queue_call_reqs => default_initializer_free_queue_call_reqs(0 downto 0),
      default_initializer_free_queue_call_acks => default_initializer_free_queue_call_acks(0 downto 0),
      default_initializer_free_queue_call_tag => default_initializer_free_queue_call_tag(0 downto 0),
      default_initializer_free_queue_return_reqs => default_initializer_free_queue_return_reqs(0 downto 0),
      default_initializer_free_queue_return_acks => default_initializer_free_queue_return_acks(0 downto 0),
      default_initializer_free_queue_return_tag => default_initializer_free_queue_return_tag(0 downto 0),
      default_initializer_free_queue_ram_call_reqs => default_initializer_free_queue_ram_call_reqs(0 downto 0),
      default_initializer_free_queue_ram_call_acks => default_initializer_free_queue_ram_call_acks(0 downto 0),
      default_initializer_free_queue_ram_call_tag => default_initializer_free_queue_ram_call_tag(0 downto 0),
      default_initializer_free_queue_ram_return_reqs => default_initializer_free_queue_ram_return_reqs(0 downto 0),
      default_initializer_free_queue_ram_return_acks => default_initializer_free_queue_ram_return_acks(0 downto 0),
      default_initializer_free_queue_ram_return_tag => default_initializer_free_queue_ram_return_tag(0 downto 0),
      default_initializer_xx_xstr_call_reqs => default_initializer_xx_xstr_call_reqs(0 downto 0),
      default_initializer_xx_xstr_call_acks => default_initializer_xx_xstr_call_acks(0 downto 0),
      default_initializer_xx_xstr_call_tag => default_initializer_xx_xstr_call_tag(0 downto 0),
      default_initializer_xx_xstr_return_reqs => default_initializer_xx_xstr_return_reqs(0 downto 0),
      default_initializer_xx_xstr_return_acks => default_initializer_xx_xstr_return_acks(0 downto 0),
      default_initializer_xx_xstr_return_tag => default_initializer_xx_xstr_return_tag(0 downto 0),
      default_initializer_xx_xstr1_call_reqs => default_initializer_xx_xstr1_call_reqs(0 downto 0),
      default_initializer_xx_xstr1_call_acks => default_initializer_xx_xstr1_call_acks(0 downto 0),
      default_initializer_xx_xstr1_call_tag => default_initializer_xx_xstr1_call_tag(0 downto 0),
      default_initializer_xx_xstr1_return_reqs => default_initializer_xx_xstr1_return_reqs(0 downto 0),
      default_initializer_xx_xstr1_return_acks => default_initializer_xx_xstr1_return_acks(0 downto 0),
      default_initializer_xx_xstr1_return_tag => default_initializer_xx_xstr1_return_tag(0 downto 0),
      default_initializer_xx_xstr2_call_reqs => default_initializer_xx_xstr2_call_reqs(0 downto 0),
      default_initializer_xx_xstr2_call_acks => default_initializer_xx_xstr2_call_acks(0 downto 0),
      default_initializer_xx_xstr2_call_tag => default_initializer_xx_xstr2_call_tag(0 downto 0),
      default_initializer_xx_xstr2_return_reqs => default_initializer_xx_xstr2_return_reqs(0 downto 0),
      default_initializer_xx_xstr2_return_acks => default_initializer_xx_xstr2_return_acks(0 downto 0),
      default_initializer_xx_xstr2_return_tag => default_initializer_xx_xstr2_return_tag(0 downto 0),
      default_initializer_xx_xstr3_call_reqs => default_initializer_xx_xstr3_call_reqs(0 downto 0),
      default_initializer_xx_xstr3_call_acks => default_initializer_xx_xstr3_call_acks(0 downto 0),
      default_initializer_xx_xstr3_call_tag => default_initializer_xx_xstr3_call_tag(0 downto 0),
      default_initializer_xx_xstr3_return_reqs => default_initializer_xx_xstr3_return_reqs(0 downto 0),
      default_initializer_xx_xstr3_return_acks => default_initializer_xx_xstr3_return_acks(0 downto 0),
      default_initializer_xx_xstr3_return_tag => default_initializer_xx_xstr3_return_tag(0 downto 0),
      default_initializer_xx_xstr4_call_reqs => default_initializer_xx_xstr4_call_reqs(0 downto 0),
      default_initializer_xx_xstr4_call_acks => default_initializer_xx_xstr4_call_acks(0 downto 0),
      default_initializer_xx_xstr4_call_tag => default_initializer_xx_xstr4_call_tag(0 downto 0),
      default_initializer_xx_xstr4_return_reqs => default_initializer_xx_xstr4_return_reqs(0 downto 0),
      default_initializer_xx_xstr4_return_acks => default_initializer_xx_xstr4_return_acks(0 downto 0),
      default_initializer_xx_xstr4_return_tag => default_initializer_xx_xstr4_return_tag(0 downto 0),
      default_initializer_xx_xstr5_call_reqs => default_initializer_xx_xstr5_call_reqs(0 downto 0),
      default_initializer_xx_xstr5_call_acks => default_initializer_xx_xstr5_call_acks(0 downto 0),
      default_initializer_xx_xstr5_call_tag => default_initializer_xx_xstr5_call_tag(0 downto 0),
      default_initializer_xx_xstr5_return_reqs => default_initializer_xx_xstr5_return_reqs(0 downto 0),
      default_initializer_xx_xstr5_return_acks => default_initializer_xx_xstr5_return_acks(0 downto 0),
      default_initializer_xx_xstr5_return_tag => default_initializer_xx_xstr5_return_tag(0 downto 0),
      default_initializer_xx_xstr6_call_reqs => default_initializer_xx_xstr6_call_reqs(0 downto 0),
      default_initializer_xx_xstr6_call_acks => default_initializer_xx_xstr6_call_acks(0 downto 0),
      default_initializer_xx_xstr6_call_tag => default_initializer_xx_xstr6_call_tag(0 downto 0),
      default_initializer_xx_xstr6_return_reqs => default_initializer_xx_xstr6_return_reqs(0 downto 0),
      default_initializer_xx_xstr6_return_acks => default_initializer_xx_xstr6_return_acks(0 downto 0),
      default_initializer_xx_xstr6_return_tag => default_initializer_xx_xstr6_return_tag(0 downto 0),
      default_initializer_xx_xstr7_call_reqs => default_initializer_xx_xstr7_call_reqs(0 downto 0),
      default_initializer_xx_xstr7_call_acks => default_initializer_xx_xstr7_call_acks(0 downto 0),
      default_initializer_xx_xstr7_call_tag => default_initializer_xx_xstr7_call_tag(0 downto 0),
      default_initializer_xx_xstr7_return_reqs => default_initializer_xx_xstr7_return_reqs(0 downto 0),
      default_initializer_xx_xstr7_return_acks => default_initializer_xx_xstr7_return_acks(0 downto 0),
      default_initializer_xx_xstr7_return_tag => default_initializer_xx_xstr7_return_tag(0 downto 0),
      default_initializer_xx_xstr8_call_reqs => default_initializer_xx_xstr8_call_reqs(0 downto 0),
      default_initializer_xx_xstr8_call_acks => default_initializer_xx_xstr8_call_acks(0 downto 0),
      default_initializer_xx_xstr8_call_tag => default_initializer_xx_xstr8_call_tag(0 downto 0),
      default_initializer_xx_xstr8_return_reqs => default_initializer_xx_xstr8_return_reqs(0 downto 0),
      default_initializer_xx_xstr8_return_acks => default_initializer_xx_xstr8_return_acks(0 downto 0),
      default_initializer_xx_xstr8_return_tag => default_initializer_xx_xstr8_return_tag(0 downto 0),
      tag_in => global_storage_initializer_x_tag_in,
      tag_out => global_storage_initializer_x_tag_out-- 
    ); -- 
  -- module wrapper_input
  wrapper_input_instance:wrapper_input-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_input_start_req,
      start_ack => wrapper_input_start_ack,
      fin_req => wrapper_input_fin_req,
      fin_ack => wrapper_input_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(7 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(7 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(87 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(15 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(7 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(7 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(15 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(3 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(7 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      free_queue_ack_pipe_read_req => free_queue_ack_pipe_read_req(0 downto 0),
      free_queue_ack_pipe_read_ack => free_queue_ack_pipe_read_ack(0 downto 0),
      free_queue_ack_pipe_read_data => free_queue_ack_pipe_read_data(7 downto 0),
      free_queue_get_pipe_read_req => free_queue_get_pipe_read_req(0 downto 0),
      free_queue_get_pipe_read_ack => free_queue_get_pipe_read_ack(0 downto 0),
      free_queue_get_pipe_read_data => free_queue_get_pipe_read_data(31 downto 0),
      in_ctrl_pipe_read_req => in_ctrl_pipe_read_req(0 downto 0),
      in_ctrl_pipe_read_ack => in_ctrl_pipe_read_ack(0 downto 0),
      in_ctrl_pipe_read_data => in_ctrl_pipe_read_data(7 downto 0),
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(1 downto 1),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(1 downto 1),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(15 downto 8),
      midpipe_pipe_write_req => midpipe_pipe_write_req(0 downto 0),
      midpipe_pipe_write_ack => midpipe_pipe_write_ack(0 downto 0),
      midpipe_pipe_write_data => midpipe_pipe_write_data(31 downto 0),
      tag_in => wrapper_input_tag_in,
      tag_out => wrapper_input_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_input_tag_in <= (others => '0');
  wrapper_input_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_input_start_req, start_ack => wrapper_input_start_ack,  fin_req => wrapper_input_fin_req,  fin_ack => wrapper_input_fin_ack);
  -- module wrapper_output
  wrapper_output_instance:wrapper_output-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_output_start_req,
      start_ack => wrapper_output_start_ack,
      fin_req => wrapper_output_fin_req,
      fin_ack => wrapper_output_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(7 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(7 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(87 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(15 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(7 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(7 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(15 downto 0),
      midpipe_pipe_read_req => midpipe_pipe_read_req(0 downto 0),
      midpipe_pipe_read_ack => midpipe_pipe_read_ack(0 downto 0),
      midpipe_pipe_read_data => midpipe_pipe_read_data(31 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(0 downto 0),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(0 downto 0),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(7 downto 0),
      free_queue_put_pipe_write_req => free_queue_put_pipe_write_req(0 downto 0),
      free_queue_put_pipe_write_ack => free_queue_put_pipe_write_ack(0 downto 0),
      free_queue_put_pipe_write_data => free_queue_put_pipe_write_data(31 downto 0),
      out_ctrl_pipe_write_req => out_ctrl_pipe_write_req(0 downto 0),
      out_ctrl_pipe_write_ack => out_ctrl_pipe_write_ack(0 downto 0),
      out_ctrl_pipe_write_data => out_ctrl_pipe_write_data(7 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(63 downto 0),
      tag_in => wrapper_output_tag_in,
      tag_out => wrapper_output_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_output_tag_in <= (others => '0');
  wrapper_output_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_output_start_req, start_ack => wrapper_output_start_ack,  fin_req => wrapper_output_fin_req,  fin_ack => wrapper_output_fin_ack);
  free_queue_ack_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_ack_pipe_read_req,
      read_ack => free_queue_ack_pipe_read_ack,
      read_data => free_queue_ack_pipe_read_data,
      write_req => free_queue_ack_pipe_write_req,
      write_ack => free_queue_ack_pipe_write_ack,
      write_data => free_queue_ack_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_get_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_get_pipe_read_req,
      read_ack => free_queue_get_pipe_read_ack,
      read_data => free_queue_get_pipe_read_data,
      write_req => free_queue_get_pipe_write_req,
      write_ack => free_queue_get_pipe_write_ack,
      write_data => free_queue_get_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_put_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_put_pipe_read_req,
      read_ack => free_queue_put_pipe_read_ack,
      read_data => free_queue_put_pipe_read_data,
      write_req => free_queue_put_pipe_write_req,
      write_ack => free_queue_put_pipe_write_ack,
      write_data => free_queue_put_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_request_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_request_pipe_read_req,
      read_ack => free_queue_request_pipe_read_ack,
      read_data => free_queue_request_pipe_read_data,
      write_req => free_queue_request_pipe_write_req,
      write_ack => free_queue_request_pipe_write_ack,
      write_data => free_queue_request_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => in_ctrl_pipe_read_req,
      read_ack => in_ctrl_pipe_read_ack,
      read_data => in_ctrl_pipe_read_data,
      write_req => in_ctrl_pipe_write_req,
      write_ack => in_ctrl_pipe_write_ack,
      write_data => in_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  midpipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => midpipe_pipe_read_req,
      read_ack => midpipe_pipe_read_ack,
      read_data => midpipe_pipe_read_data,
      write_req => midpipe_pipe_write_req,
      write_ack => midpipe_pipe_write_ack,
      write_data => midpipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => out_ctrl_pipe_read_req,
      read_ack => out_ctrl_pipe_read_ack,
      read_data => out_ctrl_pipe_read_data,
      write_req => out_ctrl_pipe_write_req,
      write_ack => out_ctrl_pipe_write_ack,
      write_data => out_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: memory_subsystem -- 
    generic map(-- 
      num_loads => 8,
      num_stores => 9,
      addr_width => 11,
      data_width => 8,
      tag_width => 2,
      number_of_banks => 4,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 2,
      addr_width => 4,
      data_width => 8,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_10: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_10_sr_addr,
      sr_data_in => memory_space_10_sr_data,
      sr_req_in => memory_space_10_sr_req,
      sr_ack_out => memory_space_10_sr_ack,
      sr_tag_in => memory_space_10_sr_tag,
      sc_req_in=> memory_space_10_sc_req,
      sc_ack_out => memory_space_10_sc_ack,
      sc_tag_out => memory_space_10_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_11: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_11_sr_addr,
      sr_data_in => memory_space_11_sr_data,
      sr_req_in => memory_space_11_sr_req,
      sr_ack_out => memory_space_11_sr_ack,
      sr_tag_in => memory_space_11_sr_tag,
      sc_req_in=> memory_space_11_sc_req,
      sc_ack_out => memory_space_11_sc_ack,
      sc_tag_out => memory_space_11_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_2: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 5,
      addr_width => 3,
      data_width => 8,
      tag_width => 2,
      num_registers => 4) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_3: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 5,
      data_width => 8,
      tag_width => 5
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_4: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_5: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_6: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_7: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_8: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_9: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 4
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
