------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai, Ch. V. Kalyani
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
--------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.types.all;
use ahir.utilities.all;

package mem_ASIC_components is

  component SZKA65_32X32X1CM2 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      DO8 : out std_logic;
      DO9 : out std_logic;
      DO10 : out std_logic;
      DO11 : out std_logic;
      DO12 : out std_logic;
      DO13 : out std_logic;
      DO14 : out std_logic;
      DO15 : out std_logic;
      DO16 : out std_logic;
      DO17 : out std_logic;
      DO18 : out std_logic;
      DO19 : out std_logic;
      DO20 : out std_logic;
      DO21 : out std_logic;
      DO22 : out std_logic;
      DO23 : out std_logic;
      DO24 : out std_logic;
      DO25 : out std_logic;
      DO26 : out std_logic;
      DO27 : out std_logic;
      DO28 : out std_logic;
      DO29 : out std_logic;
      DO30 : out std_logic;
      DO31 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      DI8 : in std_logic;
      DI9 : in std_logic;
      DI10 : in std_logic;
      DI11 : in std_logic;
      DI12 : in std_logic;
      DI13 : in std_logic;
      DI14 : in std_logic;
      DI15 : in std_logic;
      DI16 : in std_logic;
      DI17 : in std_logic;
      DI18 : in std_logic;
      DI19 : in std_logic;
      DI20 : in std_logic;
      DI21 : in std_logic;
      DI22 : in std_logic;
      DI23 : in std_logic;
      DI24 : in std_logic;
      DI25 : in std_logic;
      DI26 : in std_logic;
      DI27 : in std_logic;
      DI28 : in std_logic;
      DI29 : in std_logic;
      DI30 : in std_logic;
      DI31 : in std_logic;
      B0 : in std_logic;
      B1 : in std_logic;
      B2 : in std_logic;
      B3 : in std_logic;
      B4 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0, DVS1, DVS2:   IN   std_logic;
      CKA, CKB   :   IN   std_logic;
      CSAN, CSBN  :   IN   std_logic
);
  end component;
  component SZKA65_64X32X1CM2 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      DO8 : out std_logic;
      DO9 : out std_logic;
      DO10 : out std_logic;
      DO11 : out std_logic;
      DO12 : out std_logic;
      DO13 : out std_logic;
      DO14 : out std_logic;
      DO15 : out std_logic;
      DO16 : out std_logic;
      DO17 : out std_logic;
      DO18 : out std_logic;
      DO19 : out std_logic;
      DO20 : out std_logic;
      DO21 : out std_logic;
      DO22 : out std_logic;
      DO23 : out std_logic;
      DO24 : out std_logic;
      DO25 : out std_logic;
      DO26 : out std_logic;
      DO27 : out std_logic;
      DO28 : out std_logic;
      DO29 : out std_logic;
      DO30 : out std_logic;
      DO31 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      DI8 : in std_logic;
      DI9 : in std_logic;
      DI10 : in std_logic;
      DI11 : in std_logic;
      DI12 : in std_logic;
      DI13 : in std_logic;
      DI14 : in std_logic;
      DI15 : in std_logic;
      DI16 : in std_logic;
      DI17 : in std_logic;
      DI18 : in std_logic;
      DI19 : in std_logic;
      DI20 : in std_logic;
      DI21 : in std_logic;
      DI22 : in std_logic;
      DI23 : in std_logic;
      DI24 : in std_logic;
      DI25 : in std_logic;
      DI26 : in std_logic;
      DI27 : in std_logic;
      DI28 : in std_logic;
      DI29 : in std_logic;
      DI30 : in std_logic;
      DI31 : in std_logic;
      B0 : in std_logic;
      B1 : in std_logic;
      B2 : in std_logic;
      B3 : in std_logic;
      B4 : in std_logic;
      B5 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0, DVS1, DVS2:   IN   std_logic;
      CKA, CKB   :   IN   std_logic;
      CSAN, CSBN  :   IN   std_logic
);
  end component;
  component SHKA65_16X30X1CM4 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      DO8 : out std_logic;
      DO9 : out std_logic;
      DO10 : out std_logic;
      DO11 : out std_logic;
      DO12 : out std_logic;
      DO13 : out std_logic;
      DO14 : out std_logic;
      DO15 : out std_logic;
      DO16 : out std_logic;
      DO17 : out std_logic;
      DO18 : out std_logic;
      DO19 : out std_logic;
      DO20 : out std_logic;
      DO21 : out std_logic;
      DO22 : out std_logic;
      DO23 : out std_logic;
      DO24 : out std_logic;
      DO25 : out std_logic;
      DO26 : out std_logic;
      DO27 : out std_logic;
      DO28 : out std_logic;
      DO29 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      DI8 : in std_logic;
      DI9 : in std_logic;
      DI10 : in std_logic;
      DI11 : in std_logic;
      DI12 : in std_logic;
      DI13 : in std_logic;
      DI14 : in std_logic;
      DI15 : in std_logic;
      DI16 : in std_logic;
      DI17 : in std_logic;
      DI18 : in std_logic;
      DI19 : in std_logic;
      DI20 : in std_logic;
      DI21 : in std_logic;
      DI22 : in std_logic;
      DI23 : in std_logic;
      DI24 : in std_logic;
      DI25 : in std_logic;
      DI26 : in std_logic;
      DI27 : in std_logic;
      DI28 : in std_logic;
      DI29 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0,DVS1,DVS2:   IN   std_logic;
      CK   :   IN   std_logic;
      CSB  :   IN   std_logic
);
  end component;
  component SHKA65_32X32X1CM4 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      DO8 : out std_logic;
      DO9 : out std_logic;
      DO10 : out std_logic;
      DO11 : out std_logic;
      DO12 : out std_logic;
      DO13 : out std_logic;
      DO14 : out std_logic;
      DO15 : out std_logic;
      DO16 : out std_logic;
      DO17 : out std_logic;
      DO18 : out std_logic;
      DO19 : out std_logic;
      DO20 : out std_logic;
      DO21 : out std_logic;
      DO22 : out std_logic;
      DO23 : out std_logic;
      DO24 : out std_logic;
      DO25 : out std_logic;
      DO26 : out std_logic;
      DO27 : out std_logic;
      DO28 : out std_logic;
      DO29 : out std_logic;
      DO30 : out std_logic;
      DO31 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      DI8 : in std_logic;
      DI9 : in std_logic;
      DI10 : in std_logic;
      DI11 : in std_logic;
      DI12 : in std_logic;
      DI13 : in std_logic;
      DI14 : in std_logic;
      DI15 : in std_logic;
      DI16 : in std_logic;
      DI17 : in std_logic;
      DI18 : in std_logic;
      DI19 : in std_logic;
      DI20 : in std_logic;
      DI21 : in std_logic;
      DI22 : in std_logic;
      DI23 : in std_logic;
      DI24 : in std_logic;
      DI25 : in std_logic;
      DI26 : in std_logic;
      DI27 : in std_logic;
      DI28 : in std_logic;
      DI29 : in std_logic;
      DI30 : in std_logic;
      DI31 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0,DVS1,DVS2:   IN   std_logic;
      CK   :   IN   std_logic;
      CSB  :   IN   std_logic
);
  end component;
  component SHKA65_64X23X1CM4 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      DO8 : out std_logic;
      DO9 : out std_logic;
      DO10 : out std_logic;
      DO11 : out std_logic;
      DO12 : out std_logic;
      DO13 : out std_logic;
      DO14 : out std_logic;
      DO15 : out std_logic;
      DO16 : out std_logic;
      DO17 : out std_logic;
      DO18 : out std_logic;
      DO19 : out std_logic;
      DO20 : out std_logic;
      DO21 : out std_logic;
      DO22 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      DI8 : in std_logic;
      DI9 : in std_logic;
      DI10 : in std_logic;
      DI11 : in std_logic;
      DI12 : in std_logic;
      DI13 : in std_logic;
      DI14 : in std_logic;
      DI15 : in std_logic;
      DI16 : in std_logic;
      DI17 : in std_logic;
      DI18 : in std_logic;
      DI19 : in std_logic;
      DI20 : in std_logic;
      DI21 : in std_logic;
      DI22 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0,DVS1,DVS2:   IN   std_logic;
      CK   :   IN   std_logic;
      CSB  :   IN   std_logic
);
  end component;
  component SHKA65_512X8X1CM4 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      A6 : in std_logic;
      A7 : in std_logic;
      A8 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0,DVS1,DVS2:   IN   std_logic;
      CK   :   IN   std_logic;
      CSB  :   IN   std_logic
);
  end component;
  component SHKA65_512X64X1CM4 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      DO8 : out std_logic;
      DO9 : out std_logic;
      DO10 : out std_logic;
      DO11 : out std_logic;
      DO12 : out std_logic;
      DO13 : out std_logic;
      DO14 : out std_logic;
      DO15 : out std_logic;
      DO16 : out std_logic;
      DO17 : out std_logic;
      DO18 : out std_logic;
      DO19 : out std_logic;
      DO20 : out std_logic;
      DO21 : out std_logic;
      DO22 : out std_logic;
      DO23 : out std_logic;
      DO24 : out std_logic;
      DO25 : out std_logic;
      DO26 : out std_logic;
      DO27 : out std_logic;
      DO28 : out std_logic;
      DO29 : out std_logic;
      DO30 : out std_logic;
      DO31 : out std_logic;
      DO32 : out std_logic;
      DO33 : out std_logic;
      DO34 : out std_logic;
      DO35 : out std_logic;
      DO36 : out std_logic;
      DO37 : out std_logic;
      DO38 : out std_logic;
      DO39 : out std_logic;
      DO40 : out std_logic;
      DO41 : out std_logic;
      DO42 : out std_logic;
      DO43 : out std_logic;
      DO44 : out std_logic;
      DO45 : out std_logic;
      DO46 : out std_logic;
      DO47 : out std_logic;
      DO48 : out std_logic;
      DO49 : out std_logic;
      DO50 : out std_logic;
      DO51 : out std_logic;
      DO52 : out std_logic;
      DO53 : out std_logic;
      DO54 : out std_logic;
      DO55 : out std_logic;
      DO56 : out std_logic;
      DO57 : out std_logic;
      DO58 : out std_logic;
      DO59 : out std_logic;
      DO60 : out std_logic;
      DO61 : out std_logic;
      DO62 : out std_logic;
      DO63 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      A6 : in std_logic;
      A7 : in std_logic;
      A8 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      DI8 : in std_logic;
      DI9 : in std_logic;
      DI10 : in std_logic;
      DI11 : in std_logic;
      DI12 : in std_logic;
      DI13 : in std_logic;
      DI14 : in std_logic;
      DI15 : in std_logic;
      DI16 : in std_logic;
      DI17 : in std_logic;
      DI18 : in std_logic;
      DI19 : in std_logic;
      DI20 : in std_logic;
      DI21 : in std_logic;
      DI22 : in std_logic;
      DI23 : in std_logic;
      DI24 : in std_logic;
      DI25 : in std_logic;
      DI26 : in std_logic;
      DI27 : in std_logic;
      DI28 : in std_logic;
      DI29 : in std_logic;
      DI30 : in std_logic;
      DI31 : in std_logic;
      DI32 : in std_logic;
      DI33 : in std_logic;
      DI34 : in std_logic;
      DI35 : in std_logic;
      DI36 : in std_logic;
      DI37 : in std_logic;
      DI38 : in std_logic;
      DI39 : in std_logic;
      DI40 : in std_logic;
      DI41 : in std_logic;
      DI42 : in std_logic;
      DI43 : in std_logic;
      DI44 : in std_logic;
      DI45 : in std_logic;
      DI46 : in std_logic;
      DI47 : in std_logic;
      DI48 : in std_logic;
      DI49 : in std_logic;
      DI50 : in std_logic;
      DI51 : in std_logic;
      DI52 : in std_logic;
      DI53 : in std_logic;
      DI54 : in std_logic;
      DI55 : in std_logic;
      DI56 : in std_logic;
      DI57 : in std_logic;
      DI58 : in std_logic;
      DI59 : in std_logic;
      DI60 : in std_logic;
      DI61 : in std_logic;
      DI62 : in std_logic;
      DI63 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0,DVS1,DVS2:   IN   std_logic;
      CK   :   IN   std_logic;
      CSB  :   IN   std_logic
);
  end component;
  component SHKA65_4096X8X1CM4 is
   port(       DO0 : out std_logic;
      DO1 : out std_logic;
      DO2 : out std_logic;
      DO3 : out std_logic;
      DO4 : out std_logic;
      DO5 : out std_logic;
      DO6 : out std_logic;
      DO7 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      A6 : in std_logic;
      A7 : in std_logic;
      A8 : in std_logic;
      A9 : in std_logic;
      A10 : in std_logic;
      A11 : in std_logic;
      DI0 : in std_logic;
      DI1 : in std_logic;
      DI2 : in std_logic;
      DI3 : in std_logic;
      DI4 : in std_logic;
      DI5 : in std_logic;
      DI6 : in std_logic;
      DI7 : in std_logic;
      WEB  :   IN   std_logic;
      DVSE :   IN   std_logic;
      DVS0,DVS1,DVS2:   IN   std_logic;
      CK   :   IN   std_logic;
      CSB  :   IN   std_logic
);
  end component;
  component SJKA65_32X32X1CM4 is
   port(       DOA0 : out std_logic;
      DOA1 : out std_logic;
      DOA2 : out std_logic;
      DOA3 : out std_logic;
      DOA4 : out std_logic;
      DOA5 : out std_logic;
      DOA6 : out std_logic;
      DOA7 : out std_logic;
      DOA8 : out std_logic;
      DOA9 : out std_logic;
      DOA10 : out std_logic;
      DOA11 : out std_logic;
      DOA12 : out std_logic;
      DOA13 : out std_logic;
      DOA14 : out std_logic;
      DOA15 : out std_logic;
      DOA16 : out std_logic;
      DOA17 : out std_logic;
      DOA18 : out std_logic;
      DOA19 : out std_logic;
      DOA20 : out std_logic;
      DOA21 : out std_logic;
      DOA22 : out std_logic;
      DOA23 : out std_logic;
      DOA24 : out std_logic;
      DOA25 : out std_logic;
      DOA26 : out std_logic;
      DOA27 : out std_logic;
      DOA28 : out std_logic;
      DOA29 : out std_logic;
      DOA30 : out std_logic;
      DOA31 : out std_logic;
      DOB0 : out std_logic;
      DOB1 : out std_logic;
      DOB2 : out std_logic;
      DOB3 : out std_logic;
      DOB4 : out std_logic;
      DOB5 : out std_logic;
      DOB6 : out std_logic;
      DOB7 : out std_logic;
      DOB8 : out std_logic;
      DOB9 : out std_logic;
      DOB10 : out std_logic;
      DOB11 : out std_logic;
      DOB12 : out std_logic;
      DOB13 : out std_logic;
      DOB14 : out std_logic;
      DOB15 : out std_logic;
      DOB16 : out std_logic;
      DOB17 : out std_logic;
      DOB18 : out std_logic;
      DOB19 : out std_logic;
      DOB20 : out std_logic;
      DOB21 : out std_logic;
      DOB22 : out std_logic;
      DOB23 : out std_logic;
      DOB24 : out std_logic;
      DOB25 : out std_logic;
      DOB26 : out std_logic;
      DOB27 : out std_logic;
      DOB28 : out std_logic;
      DOB29 : out std_logic;
      DOB30 : out std_logic;
      DOB31 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      B0 : in std_logic;
      B1 : in std_logic;
      B2 : in std_logic;
      B3 : in std_logic;
      B4 : in std_logic;
      DIA0 : in std_logic;
      DIA1 : in std_logic;
      DIA2 : in std_logic;
      DIA3 : in std_logic;
      DIA4 : in std_logic;
      DIA5 : in std_logic;
      DIA6 : in std_logic;
      DIA7 : in std_logic;
      DIA8 : in std_logic;
      DIA9 : in std_logic;
      DIA10 : in std_logic;
      DIA11 : in std_logic;
      DIA12 : in std_logic;
      DIA13 : in std_logic;
      DIA14 : in std_logic;
      DIA15 : in std_logic;
      DIA16 : in std_logic;
      DIA17 : in std_logic;
      DIA18 : in std_logic;
      DIA19 : in std_logic;
      DIA20 : in std_logic;
      DIA21 : in std_logic;
      DIA22 : in std_logic;
      DIA23 : in std_logic;
      DIA24 : in std_logic;
      DIA25 : in std_logic;
      DIA26 : in std_logic;
      DIA27 : in std_logic;
      DIA28 : in std_logic;
      DIA29 : in std_logic;
      DIA30 : in std_logic;
      DIA31 : in std_logic;
      DIB0 : in std_logic;
      DIB1 : in std_logic;
      DIB2 : in std_logic;
      DIB3 : in std_logic;
      DIB4 : in std_logic;
      DIB5 : in std_logic;
      DIB6 : in std_logic;
      DIB7 : in std_logic;
      DIB8 : in std_logic;
      DIB9 : in std_logic;
      DIB10 : in std_logic;
      DIB11 : in std_logic;
      DIB12 : in std_logic;
      DIB13 : in std_logic;
      DIB14 : in std_logic;
      DIB15 : in std_logic;
      DIB16 : in std_logic;
      DIB17 : in std_logic;
      DIB18 : in std_logic;
      DIB19 : in std_logic;
      DIB20 : in std_logic;
      DIB21 : in std_logic;
      DIB22 : in std_logic;
      DIB23 : in std_logic;
      DIB24 : in std_logic;
      DIB25 : in std_logic;
      DIB26 : in std_logic;
      DIB27 : in std_logic;
      DIB28 : in std_logic;
      DIB29 : in std_logic;
      DIB30 : in std_logic;
      DIB31 : in std_logic;
     WEAN                          :   IN   std_logic;
     WEBN                          :   IN   std_logic;
     DVSE                          :   IN   std_logic;
     DVS0, DVS1, DVS2, DVS3        :   IN   std_logic;
     CKA                           :   IN   std_logic;
     CKB                           :   IN   std_logic;
     CSAN                          :   IN   std_logic;
     CSBN                          :   IN   std_logic
);
  end component;
  component SJKA65_64X32X1CM4 is
   port(       DOA0 : out std_logic;
      DOA1 : out std_logic;
      DOA2 : out std_logic;
      DOA3 : out std_logic;
      DOA4 : out std_logic;
      DOA5 : out std_logic;
      DOA6 : out std_logic;
      DOA7 : out std_logic;
      DOA8 : out std_logic;
      DOA9 : out std_logic;
      DOA10 : out std_logic;
      DOA11 : out std_logic;
      DOA12 : out std_logic;
      DOA13 : out std_logic;
      DOA14 : out std_logic;
      DOA15 : out std_logic;
      DOA16 : out std_logic;
      DOA17 : out std_logic;
      DOA18 : out std_logic;
      DOA19 : out std_logic;
      DOA20 : out std_logic;
      DOA21 : out std_logic;
      DOA22 : out std_logic;
      DOA23 : out std_logic;
      DOA24 : out std_logic;
      DOA25 : out std_logic;
      DOA26 : out std_logic;
      DOA27 : out std_logic;
      DOA28 : out std_logic;
      DOA29 : out std_logic;
      DOA30 : out std_logic;
      DOA31 : out std_logic;
      DOB0 : out std_logic;
      DOB1 : out std_logic;
      DOB2 : out std_logic;
      DOB3 : out std_logic;
      DOB4 : out std_logic;
      DOB5 : out std_logic;
      DOB6 : out std_logic;
      DOB7 : out std_logic;
      DOB8 : out std_logic;
      DOB9 : out std_logic;
      DOB10 : out std_logic;
      DOB11 : out std_logic;
      DOB12 : out std_logic;
      DOB13 : out std_logic;
      DOB14 : out std_logic;
      DOB15 : out std_logic;
      DOB16 : out std_logic;
      DOB17 : out std_logic;
      DOB18 : out std_logic;
      DOB19 : out std_logic;
      DOB20 : out std_logic;
      DOB21 : out std_logic;
      DOB22 : out std_logic;
      DOB23 : out std_logic;
      DOB24 : out std_logic;
      DOB25 : out std_logic;
      DOB26 : out std_logic;
      DOB27 : out std_logic;
      DOB28 : out std_logic;
      DOB29 : out std_logic;
      DOB30 : out std_logic;
      DOB31 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      B0 : in std_logic;
      B1 : in std_logic;
      B2 : in std_logic;
      B3 : in std_logic;
      B4 : in std_logic;
      B5 : in std_logic;
      DIA0 : in std_logic;
      DIA1 : in std_logic;
      DIA2 : in std_logic;
      DIA3 : in std_logic;
      DIA4 : in std_logic;
      DIA5 : in std_logic;
      DIA6 : in std_logic;
      DIA7 : in std_logic;
      DIA8 : in std_logic;
      DIA9 : in std_logic;
      DIA10 : in std_logic;
      DIA11 : in std_logic;
      DIA12 : in std_logic;
      DIA13 : in std_logic;
      DIA14 : in std_logic;
      DIA15 : in std_logic;
      DIA16 : in std_logic;
      DIA17 : in std_logic;
      DIA18 : in std_logic;
      DIA19 : in std_logic;
      DIA20 : in std_logic;
      DIA21 : in std_logic;
      DIA22 : in std_logic;
      DIA23 : in std_logic;
      DIA24 : in std_logic;
      DIA25 : in std_logic;
      DIA26 : in std_logic;
      DIA27 : in std_logic;
      DIA28 : in std_logic;
      DIA29 : in std_logic;
      DIA30 : in std_logic;
      DIA31 : in std_logic;
      DIB0 : in std_logic;
      DIB1 : in std_logic;
      DIB2 : in std_logic;
      DIB3 : in std_logic;
      DIB4 : in std_logic;
      DIB5 : in std_logic;
      DIB6 : in std_logic;
      DIB7 : in std_logic;
      DIB8 : in std_logic;
      DIB9 : in std_logic;
      DIB10 : in std_logic;
      DIB11 : in std_logic;
      DIB12 : in std_logic;
      DIB13 : in std_logic;
      DIB14 : in std_logic;
      DIB15 : in std_logic;
      DIB16 : in std_logic;
      DIB17 : in std_logic;
      DIB18 : in std_logic;
      DIB19 : in std_logic;
      DIB20 : in std_logic;
      DIB21 : in std_logic;
      DIB22 : in std_logic;
      DIB23 : in std_logic;
      DIB24 : in std_logic;
      DIB25 : in std_logic;
      DIB26 : in std_logic;
      DIB27 : in std_logic;
      DIB28 : in std_logic;
      DIB29 : in std_logic;
      DIB30 : in std_logic;
      DIB31 : in std_logic;
     WEAN                          :   IN   std_logic;
     WEBN                          :   IN   std_logic;
     DVSE                          :   IN   std_logic;
     DVS0, DVS1, DVS2, DVS3        :   IN   std_logic;
     CKA                           :   IN   std_logic;
     CKB                           :   IN   std_logic;
     CSAN                          :   IN   std_logic;
     CSBN                          :   IN   std_logic
);
  end component;
  component SJKA65_256X54X1CM4 is
   port(       DOA0 : out std_logic;
      DOA1 : out std_logic;
      DOA2 : out std_logic;
      DOA3 : out std_logic;
      DOA4 : out std_logic;
      DOA5 : out std_logic;
      DOA6 : out std_logic;
      DOA7 : out std_logic;
      DOA8 : out std_logic;
      DOA9 : out std_logic;
      DOA10 : out std_logic;
      DOA11 : out std_logic;
      DOA12 : out std_logic;
      DOA13 : out std_logic;
      DOA14 : out std_logic;
      DOA15 : out std_logic;
      DOA16 : out std_logic;
      DOA17 : out std_logic;
      DOA18 : out std_logic;
      DOA19 : out std_logic;
      DOA20 : out std_logic;
      DOA21 : out std_logic;
      DOA22 : out std_logic;
      DOA23 : out std_logic;
      DOA24 : out std_logic;
      DOA25 : out std_logic;
      DOA26 : out std_logic;
      DOA27 : out std_logic;
      DOA28 : out std_logic;
      DOA29 : out std_logic;
      DOA30 : out std_logic;
      DOA31 : out std_logic;
      DOA32 : out std_logic;
      DOA33 : out std_logic;
      DOA34 : out std_logic;
      DOA35 : out std_logic;
      DOA36 : out std_logic;
      DOA37 : out std_logic;
      DOA38 : out std_logic;
      DOA39 : out std_logic;
      DOA40 : out std_logic;
      DOA41 : out std_logic;
      DOA42 : out std_logic;
      DOA43 : out std_logic;
      DOA44 : out std_logic;
      DOA45 : out std_logic;
      DOA46 : out std_logic;
      DOA47 : out std_logic;
      DOA48 : out std_logic;
      DOA49 : out std_logic;
      DOA50 : out std_logic;
      DOA51 : out std_logic;
      DOA52 : out std_logic;
      DOA53 : out std_logic;
      DOB0 : out std_logic;
      DOB1 : out std_logic;
      DOB2 : out std_logic;
      DOB3 : out std_logic;
      DOB4 : out std_logic;
      DOB5 : out std_logic;
      DOB6 : out std_logic;
      DOB7 : out std_logic;
      DOB8 : out std_logic;
      DOB9 : out std_logic;
      DOB10 : out std_logic;
      DOB11 : out std_logic;
      DOB12 : out std_logic;
      DOB13 : out std_logic;
      DOB14 : out std_logic;
      DOB15 : out std_logic;
      DOB16 : out std_logic;
      DOB17 : out std_logic;
      DOB18 : out std_logic;
      DOB19 : out std_logic;
      DOB20 : out std_logic;
      DOB21 : out std_logic;
      DOB22 : out std_logic;
      DOB23 : out std_logic;
      DOB24 : out std_logic;
      DOB25 : out std_logic;
      DOB26 : out std_logic;
      DOB27 : out std_logic;
      DOB28 : out std_logic;
      DOB29 : out std_logic;
      DOB30 : out std_logic;
      DOB31 : out std_logic;
      DOB32 : out std_logic;
      DOB33 : out std_logic;
      DOB34 : out std_logic;
      DOB35 : out std_logic;
      DOB36 : out std_logic;
      DOB37 : out std_logic;
      DOB38 : out std_logic;
      DOB39 : out std_logic;
      DOB40 : out std_logic;
      DOB41 : out std_logic;
      DOB42 : out std_logic;
      DOB43 : out std_logic;
      DOB44 : out std_logic;
      DOB45 : out std_logic;
      DOB46 : out std_logic;
      DOB47 : out std_logic;
      DOB48 : out std_logic;
      DOB49 : out std_logic;
      DOB50 : out std_logic;
      DOB51 : out std_logic;
      DOB52 : out std_logic;
      DOB53 : out std_logic;
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      A6 : in std_logic;
      A7 : in std_logic;
      B0 : in std_logic;
      B1 : in std_logic;
      B2 : in std_logic;
      B3 : in std_logic;
      B4 : in std_logic;
      B5 : in std_logic;
      B6 : in std_logic;
      B7 : in std_logic;
      DIA0 : in std_logic;
      DIA1 : in std_logic;
      DIA2 : in std_logic;
      DIA3 : in std_logic;
      DIA4 : in std_logic;
      DIA5 : in std_logic;
      DIA6 : in std_logic;
      DIA7 : in std_logic;
      DIA8 : in std_logic;
      DIA9 : in std_logic;
      DIA10 : in std_logic;
      DIA11 : in std_logic;
      DIA12 : in std_logic;
      DIA13 : in std_logic;
      DIA14 : in std_logic;
      DIA15 : in std_logic;
      DIA16 : in std_logic;
      DIA17 : in std_logic;
      DIA18 : in std_logic;
      DIA19 : in std_logic;
      DIA20 : in std_logic;
      DIA21 : in std_logic;
      DIA22 : in std_logic;
      DIA23 : in std_logic;
      DIA24 : in std_logic;
      DIA25 : in std_logic;
      DIA26 : in std_logic;
      DIA27 : in std_logic;
      DIA28 : in std_logic;
      DIA29 : in std_logic;
      DIA30 : in std_logic;
      DIA31 : in std_logic;
      DIA32 : in std_logic;
      DIA33 : in std_logic;
      DIA34 : in std_logic;
      DIA35 : in std_logic;
      DIA36 : in std_logic;
      DIA37 : in std_logic;
      DIA38 : in std_logic;
      DIA39 : in std_logic;
      DIA40 : in std_logic;
      DIA41 : in std_logic;
      DIA42 : in std_logic;
      DIA43 : in std_logic;
      DIA44 : in std_logic;
      DIA45 : in std_logic;
      DIA46 : in std_logic;
      DIA47 : in std_logic;
      DIA48 : in std_logic;
      DIA49 : in std_logic;
      DIA50 : in std_logic;
      DIA51 : in std_logic;
      DIA52 : in std_logic;
      DIA53 : in std_logic;
      DIB0 : in std_logic;
      DIB1 : in std_logic;
      DIB2 : in std_logic;
      DIB3 : in std_logic;
      DIB4 : in std_logic;
      DIB5 : in std_logic;
      DIB6 : in std_logic;
      DIB7 : in std_logic;
      DIB8 : in std_logic;
      DIB9 : in std_logic;
      DIB10 : in std_logic;
      DIB11 : in std_logic;
      DIB12 : in std_logic;
      DIB13 : in std_logic;
      DIB14 : in std_logic;
      DIB15 : in std_logic;
      DIB16 : in std_logic;
      DIB17 : in std_logic;
      DIB18 : in std_logic;
      DIB19 : in std_logic;
      DIB20 : in std_logic;
      DIB21 : in std_logic;
      DIB22 : in std_logic;
      DIB23 : in std_logic;
      DIB24 : in std_logic;
      DIB25 : in std_logic;
      DIB26 : in std_logic;
      DIB27 : in std_logic;
      DIB28 : in std_logic;
      DIB29 : in std_logic;
      DIB30 : in std_logic;
      DIB31 : in std_logic;
      DIB32 : in std_logic;
      DIB33 : in std_logic;
      DIB34 : in std_logic;
      DIB35 : in std_logic;
      DIB36 : in std_logic;
      DIB37 : in std_logic;
      DIB38 : in std_logic;
      DIB39 : in std_logic;
      DIB40 : in std_logic;
      DIB41 : in std_logic;
      DIB42 : in std_logic;
      DIB43 : in std_logic;
      DIB44 : in std_logic;
      DIB45 : in std_logic;
      DIB46 : in std_logic;
      DIB47 : in std_logic;
      DIB48 : in std_logic;
      DIB49 : in std_logic;
      DIB50 : in std_logic;
      DIB51 : in std_logic;
      DIB52 : in std_logic;
      DIB53 : in std_logic;
     WEAN                          :   IN   std_logic;
     WEBN                          :   IN   std_logic;
     DVSE                          :   IN   std_logic;
     DVS0, DVS1, DVS2, DVS3        :   IN   std_logic;
     CKA                           :   IN   std_logic;
     CKB                           :   IN   std_logic;
     CSAN                          :   IN   std_logic;
     CSBN                          :   IN   std_logic
);
  end component;
end package;

