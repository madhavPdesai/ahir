-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity mmultiply is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(8 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(8 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
    in_data_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    result_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    result_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    result_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    mmultiply_base_call_reqs : out  std_logic_vector(0 downto 0);
    mmultiply_base_call_acks : in   std_logic_vector(0 downto 0);
    mmultiply_base_call_tag  :  out  std_logic_vector(0 downto 0);
    mmultiply_base_return_reqs : out  std_logic_vector(0 downto 0);
    mmultiply_base_return_acks : in   std_logic_vector(0 downto 0);
    mmultiply_base_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity mmultiply;
architecture Default of mmultiply is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal mmultiply_CP_10911_start: Boolean;
  -- links between control-path and data-path
  signal simple_obj_ref_353_inst_req_0 : boolean;
  signal binary_382_inst_req_1 : boolean;
  signal ptr_deref_356_base_resize_ack_0 : boolean;
  signal simple_obj_ref_353_inst_ack_0 : boolean;
  signal binary_369_inst_ack_1 : boolean;
  signal binary_369_inst_req_1 : boolean;
  signal array_obj_ref_430_index_sum_1_req_1 : boolean;
  signal binary_388_inst_req_1 : boolean;
  signal array_obj_ref_430_index_0_resize_ack_0 : boolean;
  signal ptr_deref_356_base_resize_req_0 : boolean;
  signal if_stmt_371_branch_ack_1 : boolean;
  signal binary_388_inst_req_0 : boolean;
  signal array_obj_ref_430_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_349_root_address_inst_req_0 : boolean;
  signal array_obj_ref_430_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_430_index_sum_1_ack_1 : boolean;
  signal ptr_deref_356_store_0_ack_0 : boolean;
  signal ptr_deref_356_store_0_req_0 : boolean;
  signal ptr_deref_356_store_0_req_1 : boolean;
  signal binary_369_inst_ack_0 : boolean;
  signal ptr_deref_356_root_address_inst_req_0 : boolean;
  signal ptr_deref_437_root_address_inst_req_0 : boolean;
  signal array_obj_ref_349_index_0_scale_req_0 : boolean;
  signal array_obj_ref_430_index_0_scale_ack_0 : boolean;
  signal binary_388_inst_ack_0 : boolean;
  signal if_stmt_390_branch_req_0 : boolean;
  signal if_stmt_371_branch_req_0 : boolean;
  signal array_obj_ref_430_offset_inst_ack_0 : boolean;
  signal binary_450_inst_ack_0 : boolean;
  signal binary_382_inst_ack_1 : boolean;
  signal array_obj_ref_430_index_0_scale_req_1 : boolean;
  signal array_obj_ref_430_offset_inst_req_0 : boolean;
  signal array_obj_ref_349_index_0_scale_ack_0 : boolean;
  signal ptr_deref_356_store_0_ack_1 : boolean;
  signal array_obj_ref_349_index_0_scale_req_1 : boolean;
  signal array_obj_ref_430_index_1_rename_req_0 : boolean;
  signal array_obj_ref_430_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_430_index_0_resize_req_0 : boolean;
  signal binary_363_inst_req_1 : boolean;
  signal array_obj_ref_349_index_0_resize_req_0 : boolean;
  signal array_obj_ref_349_index_0_resize_ack_0 : boolean;
  signal binary_363_inst_ack_1 : boolean;
  signal ptr_deref_356_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_349_index_1_resize_req_0 : boolean;
  signal binary_382_inst_req_0 : boolean;
  signal binary_382_inst_ack_0 : boolean;
  signal array_obj_ref_349_root_address_inst_ack_0 : boolean;
  signal binary_444_inst_ack_1 : boolean;
  signal binary_369_inst_req_0 : boolean;
  signal array_obj_ref_349_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_349_index_sum_1_req_1 : boolean;
  signal array_obj_ref_349_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_430_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_349_offset_inst_req_0 : boolean;
  signal array_obj_ref_349_offset_inst_ack_0 : boolean;
  signal addr_of_431_final_reg_ack_0 : boolean;
  signal phi_stmt_419_ack_0 : boolean;
  signal phi_stmt_481_ack_0 : boolean;
  signal phi_stmt_419_req_0 : boolean;
  signal binary_444_inst_req_0 : boolean;
  signal binary_463_inst_req_0 : boolean;
  signal binary_463_inst_ack_0 : boolean;
  signal binary_463_inst_req_1 : boolean;
  signal binary_463_inst_ack_1 : boolean;
  signal phi_stmt_409_req_1 : boolean;
  signal binary_469_inst_req_0 : boolean;
  signal binary_469_inst_ack_0 : boolean;
  signal ptr_deref_437_store_0_ack_1 : boolean;
  signal binary_363_inst_req_0 : boolean;
  signal array_obj_ref_349_index_0_scale_ack_1 : boolean;
  signal ptr_deref_437_root_address_inst_ack_0 : boolean;
  signal ptr_deref_437_addr_0_req_0 : boolean;
  signal ptr_deref_437_addr_0_ack_0 : boolean;
  signal ptr_deref_437_store_0_req_0 : boolean;
  signal array_obj_ref_349_index_1_resize_ack_0 : boolean;
  signal ptr_deref_356_gather_scatter_req_0 : boolean;
  signal binary_444_inst_req_1 : boolean;
  signal type_cast_412_inst_ack_0 : boolean;
  signal type_cast_412_inst_req_0 : boolean;
  signal if_stmt_390_branch_ack_0 : boolean;
  signal binary_388_inst_ack_1 : boolean;
  signal ptr_deref_437_store_0_req_1 : boolean;
  signal ptr_deref_356_addr_0_req_0 : boolean;
  signal ptr_deref_437_base_resize_ack_0 : boolean;
  signal binary_444_inst_ack_0 : boolean;
  signal ptr_deref_356_addr_0_ack_0 : boolean;
  signal array_obj_ref_430_root_address_inst_req_0 : boolean;
  signal ptr_deref_437_store_0_ack_0 : boolean;
  signal ptr_deref_356_gather_scatter_ack_0 : boolean;
  signal binary_363_inst_ack_0 : boolean;
  signal if_stmt_452_branch_req_0 : boolean;
  signal array_obj_ref_349_index_1_rename_req_0 : boolean;
  signal array_obj_ref_349_index_1_rename_ack_0 : boolean;
  signal binary_450_inst_ack_1 : boolean;
  signal addr_of_350_final_reg_req_0 : boolean;
  signal array_obj_ref_430_root_address_inst_ack_0 : boolean;
  signal if_stmt_452_branch_ack_0 : boolean;
  signal binary_450_inst_req_0 : boolean;
  signal array_obj_ref_430_index_0_scale_req_0 : boolean;
  signal ptr_deref_437_gather_scatter_req_0 : boolean;
  signal phi_stmt_409_ack_0 : boolean;
  signal if_stmt_371_branch_ack_0 : boolean;
  signal addr_of_431_final_reg_req_0 : boolean;
  signal array_obj_ref_430_index_1_resize_req_0 : boolean;
  signal if_stmt_452_branch_ack_1 : boolean;
  signal addr_of_350_final_reg_ack_0 : boolean;
  signal ptr_deref_437_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_430_index_sum_1_req_0 : boolean;
  signal ptr_deref_437_base_resize_req_0 : boolean;
  signal array_obj_ref_349_index_sum_1_req_0 : boolean;
  signal if_stmt_390_branch_ack_1 : boolean;
  signal phi_stmt_409_req_0 : boolean;
  signal simple_obj_ref_434_inst_ack_0 : boolean;
  signal simple_obj_ref_434_inst_req_0 : boolean;
  signal binary_450_inst_req_1 : boolean;
  signal phi_stmt_491_ack_0 : boolean;
  signal phi_stmt_481_req_1 : boolean;
  signal type_cast_487_inst_req_0 : boolean;
  signal type_cast_425_inst_req_0 : boolean;
  signal type_cast_425_inst_ack_0 : boolean;
  signal phi_stmt_419_req_1 : boolean;
  signal type_cast_487_inst_ack_0 : boolean;
  signal binary_469_inst_req_1 : boolean;
  signal binary_469_inst_ack_1 : boolean;
  signal if_stmt_471_branch_req_0 : boolean;
  signal if_stmt_471_branch_ack_1 : boolean;
  signal if_stmt_471_branch_ack_0 : boolean;
  signal call_stmt_478_call_req_0 : boolean;
  signal call_stmt_478_call_ack_0 : boolean;
  signal call_stmt_478_call_req_1 : boolean;
  signal call_stmt_478_call_ack_1 : boolean;
  signal array_obj_ref_502_index_0_resize_req_0 : boolean;
  signal array_obj_ref_502_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_502_index_0_scale_req_0 : boolean;
  signal array_obj_ref_502_index_0_scale_ack_0 : boolean;
  signal phi_stmt_397_ack_0 : boolean;
  signal array_obj_ref_502_index_0_scale_req_1 : boolean;
  signal array_obj_ref_502_index_0_scale_ack_1 : boolean;
  signal phi_stmt_397_req_0 : boolean;
  signal type_cast_400_inst_ack_0 : boolean;
  signal type_cast_400_inst_req_0 : boolean;
  signal phi_stmt_491_req_0 : boolean;
  signal array_obj_ref_502_index_1_resize_req_0 : boolean;
  signal array_obj_ref_502_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_502_index_1_rename_req_0 : boolean;
  signal array_obj_ref_502_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_502_index_sum_1_req_0 : boolean;
  signal array_obj_ref_502_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_502_index_sum_1_req_1 : boolean;
  signal array_obj_ref_502_index_sum_1_ack_1 : boolean;
  signal phi_stmt_397_req_1 : boolean;
  signal array_obj_ref_502_offset_inst_req_0 : boolean;
  signal array_obj_ref_502_offset_inst_ack_0 : boolean;
  signal array_obj_ref_502_root_address_inst_req_0 : boolean;
  signal array_obj_ref_502_root_address_inst_ack_0 : boolean;
  signal addr_of_503_final_reg_req_0 : boolean;
  signal addr_of_503_final_reg_ack_0 : boolean;
  signal ptr_deref_507_base_resize_req_0 : boolean;
  signal ptr_deref_507_base_resize_ack_0 : boolean;
  signal ptr_deref_507_root_address_inst_req_0 : boolean;
  signal ptr_deref_507_root_address_inst_ack_0 : boolean;
  signal ptr_deref_507_addr_0_req_0 : boolean;
  signal ptr_deref_507_addr_0_ack_0 : boolean;
  signal ptr_deref_507_load_0_req_0 : boolean;
  signal phi_stmt_338_ack_0 : boolean;
  signal ptr_deref_507_load_0_ack_0 : boolean;
  signal ptr_deref_507_load_0_req_1 : boolean;
  signal ptr_deref_507_load_0_ack_1 : boolean;
  signal phi_stmt_338_req_0 : boolean;
  signal ptr_deref_507_gather_scatter_req_0 : boolean;
  signal ptr_deref_507_gather_scatter_ack_0 : boolean;
  signal phi_stmt_491_req_1 : boolean;
  signal simple_obj_ref_509_inst_req_0 : boolean;
  signal simple_obj_ref_509_inst_ack_0 : boolean;
  signal type_cast_497_inst_ack_0 : boolean;
  signal phi_stmt_338_req_1 : boolean;
  signal type_cast_344_inst_ack_0 : boolean;
  signal type_cast_344_inst_req_0 : boolean;
  signal type_cast_497_inst_req_0 : boolean;
  signal binary_516_inst_req_0 : boolean;
  signal binary_516_inst_ack_0 : boolean;
  signal binary_516_inst_req_1 : boolean;
  signal binary_516_inst_ack_1 : boolean;
  signal phi_stmt_328_ack_0 : boolean;
  signal phi_stmt_328_req_1 : boolean;
  signal type_cast_334_inst_ack_0 : boolean;
  signal type_cast_334_inst_req_0 : boolean;
  signal binary_522_inst_req_0 : boolean;
  signal binary_522_inst_ack_0 : boolean;
  signal binary_522_inst_req_1 : boolean;
  signal binary_522_inst_ack_1 : boolean;
  signal if_stmt_524_branch_req_0 : boolean;
  signal if_stmt_524_branch_ack_1 : boolean;
  signal phi_stmt_328_req_0 : boolean;
  signal if_stmt_524_branch_ack_0 : boolean;
  signal phi_stmt_481_req_0 : boolean;
  signal binary_535_inst_req_0 : boolean;
  signal binary_535_inst_ack_0 : boolean;
  signal binary_535_inst_req_1 : boolean;
  signal binary_535_inst_ack_1 : boolean;
  signal binary_541_inst_req_0 : boolean;
  signal binary_541_inst_ack_0 : boolean;
  signal binary_541_inst_req_1 : boolean;
  signal binary_541_inst_ack_1 : boolean;
  signal if_stmt_543_branch_req_0 : boolean;
  signal if_stmt_543_branch_ack_1 : boolean;
  signal if_stmt_543_branch_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  mmultiply_CP_10911: Block -- control-path 
    signal cp_elements: BooleanArray(284 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(240);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(240), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  output  bypass 
    -- predecessors 
    -- successors 248 
    -- members (15) 
      -- 	$entry
      -- 	branch_block_stmt_323/$entry
      -- 	branch_block_stmt_323/branch_block_stmt_323__entry__
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_req
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/ack
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/req
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/$exit
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/$entry
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/$entry
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/$exit
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/$entry
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/$exit
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/$entry
      -- 	branch_block_stmt_323/bb_0_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/$exit
      -- 
    phi_stmt_328_req_11778_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => phi_stmt_328_req_0); -- 
    -- CP-element group 1 branch  place  bypass 
    -- predecessors 58 
    -- successors 59 62 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370__exit__
      -- 	branch_block_stmt_323/if_stmt_371__entry__
      -- 
    cp_elements(1) <= cp_elements(58);
    -- CP-element group 2 merge  fork  transition  place  no-bypass 
    -- predecessors 65 256 
    -- successors 70 68 
    -- members (7) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/$entry
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/simple_obj_ref_379_completed_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_trigger_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/simple_obj_ref_379_trigger_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/simple_obj_ref_379_active_
      -- 	branch_block_stmt_323/merge_stmt_377__exit__
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389__entry__
      -- 
    cp_elements(2) <= OrReduce(cp_elements(65) & cp_elements(256));
    -- CP-element group 3 merge  transition  place  output  bypass 
    -- predecessors 258 262 
    -- successors 247 
    -- members (7) 
      -- 	branch_block_stmt_323/merge_stmt_396__exit__
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/req
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/$entry
      -- 
    cp_elements(3) <= OrReduce(cp_elements(258) & cp_elements(262));
    req_11791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => type_cast_334_inst_req_0); -- 
    -- CP-element group 4 branch  place  bypass 
    -- predecessors 139 
    -- successors 140 143 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451__exit__
      -- 	branch_block_stmt_323/if_stmt_452__entry__
      -- 
    cp_elements(4) <= cp_elements(139);
    -- CP-element group 5 merge  fork  transition  place  no-bypass 
    -- predecessors 146 272 
    -- successors 149 151 
    -- members (7) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/simple_obj_ref_460_trigger_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/simple_obj_ref_460_active_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/simple_obj_ref_460_completed_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_trigger_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/$entry
      -- 	branch_block_stmt_323/merge_stmt_458__exit__
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470__entry__
      -- 
    cp_elements(5) <= OrReduce(cp_elements(146) & cp_elements(272));
    -- CP-element group 6 merge  transition  place  output  bypass 
    -- predecessors 167 274 
    -- successors 170 
    -- members (6) 
      -- 	branch_block_stmt_323/merge_stmt_477__exit__
      -- 	branch_block_stmt_323/call_stmt_478__entry__
      -- 	branch_block_stmt_323/call_stmt_478/$entry
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_trigger_
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_start/$entry
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_start/crr
      -- 
    cp_elements(6) <= OrReduce(cp_elements(167) & cp_elements(274));
    crr_11497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => call_stmt_478_call_req_0); -- 
    -- CP-element group 7 merge  fork  transition  place  no-bypass 
    -- predecessors 223 284 
    -- successors 226 228 
    -- members (7) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542__entry__
      -- 	branch_block_stmt_323/merge_stmt_530__exit__
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/$entry
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_trigger_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/simple_obj_ref_532_trigger_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/simple_obj_ref_532_active_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/simple_obj_ref_532_completed_
      -- 
    cp_elements(7) <= OrReduce(cp_elements(223) & cp_elements(284));
    -- CP-element group 8 fork  transition  bypass 
    -- predecessors 254 
    -- successors 13 9 17 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_351/$entry
      -- 
    cp_elements(8) <= cp_elements(254);
    -- CP-element group 9 transition  bypass 
    -- predecessors 8 
    -- successors 10 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_351/addr_of_350_trigger_
      -- 
    cp_elements(9) <= cp_elements(8);
    -- CP-element group 10 join  fork  transition  bypass 
    -- predecessors 23 9 
    -- successors 11 24 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_351/addr_of_350_active_
      -- 
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(23);
      predecessors(1) <= cp_elements(9);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(10)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 11 join  fork  transition  place  no-bypass 
    -- predecessors 10 25 
    -- successors 27 26 
    -- members (10) 
      -- 	branch_block_stmt_323/assign_stmt_351/addr_of_350_completed_
      -- 	branch_block_stmt_323/assign_stmt_354/simple_obj_ref_353_active_
      -- 	branch_block_stmt_323/assign_stmt_354/simple_obj_ref_353_trigger_
      -- 	branch_block_stmt_323/assign_stmt_354/$entry
      -- 	branch_block_stmt_323/assign_stmt_351/assign_stmt_351_active_
      -- 	branch_block_stmt_323/assign_stmt_351/assign_stmt_351_trigger_
      -- 	branch_block_stmt_323/assign_stmt_351/$exit
      -- 	branch_block_stmt_323/assign_stmt_351/assign_stmt_351_completed_
      -- 	branch_block_stmt_323/assign_stmt_351__exit__
      -- 	branch_block_stmt_323/assign_stmt_354__entry__
      -- 
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(10);
      predecessors(1) <= cp_elements(25);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(11)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 12 join  transition  output  bypass 
    -- predecessors 19 16 
    -- successors 20 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_indices_scaled
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/$entry
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_12 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(19);
      predecessors(1) <= cp_elements(16);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(12)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(12),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_11030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => array_obj_ref_349_index_sum_1_req_0); -- 
    -- CP-element group 13 transition  output  bypass 
    -- predecessors 8 
    -- successors 14 
    -- members (6) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_computed_0
      -- 	branch_block_stmt_323/assign_stmt_351/simple_obj_ref_347_trigger_
      -- 	branch_block_stmt_323/assign_stmt_351/simple_obj_ref_347_active_
      -- 	branch_block_stmt_323/assign_stmt_351/simple_obj_ref_347_completed_
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_0/index_resize_req
      -- 
    cp_elements(13) <= cp_elements(8);
    index_resize_req_11003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => array_obj_ref_349_index_0_resize_req_0); -- 
    -- CP-element group 14 transition  input  output  no-bypass 
    -- predecessors 13 
    -- successors 15 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resized_0
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_0/scale_rr
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_0/$entry
      -- 
    index_resize_ack_11004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_index_0_resize_ack_0, ack => cp_elements(14)); -- 
    scale_rr_11008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => array_obj_ref_349_index_0_scale_req_0); -- 
    -- CP-element group 15 transition  input  output  no-bypass 
    -- predecessors 14 
    -- successors 16 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_0/scale_ra
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_0/scale_cr
      -- 
    scale_ra_11009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_index_0_scale_ack_0, ack => cp_elements(15)); -- 
    scale_cr_11010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => array_obj_ref_349_index_0_scale_req_1); -- 
    -- CP-element group 16 transition  input  no-bypass 
    -- predecessors 15 
    -- successors 12 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_0/scale_ca
      -- 
    scale_ca_11011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_index_0_scale_ack_1, ack => cp_elements(16)); -- 
    -- CP-element group 17 transition  output  bypass 
    -- predecessors 8 
    -- successors 18 
    -- members (6) 
      -- 	branch_block_stmt_323/assign_stmt_351/simple_obj_ref_348_completed_
      -- 	branch_block_stmt_323/assign_stmt_351/simple_obj_ref_348_active_
      -- 	branch_block_stmt_323/assign_stmt_351/simple_obj_ref_348_trigger_
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_1/$entry
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_1/index_resize_req
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_computed_1
      -- 
    cp_elements(17) <= cp_elements(8);
    index_resize_req_11020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => array_obj_ref_349_index_1_resize_req_0); -- 
    -- CP-element group 18 transition  input  output  no-bypass 
    -- predecessors 17 
    -- successors 19 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resized_1
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_1/$exit
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_1/$entry
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_11021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_index_1_resize_ack_0, ack => cp_elements(18)); -- 
    scale_rename_req_11025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => array_obj_ref_349_index_1_rename_req_0); -- 
    -- CP-element group 19 transition  input  no-bypass 
    -- predecessors 18 
    -- successors 12 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_1/$exit
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_11026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_index_1_rename_ack_0, ack => cp_elements(19)); -- 
    -- CP-element group 20 transition  input  output  no-bypass 
    -- predecessors 12 
    -- successors 21 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_11031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_index_sum_1_ack_0, ack => cp_elements(20)); -- 
    partial_sum_1_cr_11032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => array_obj_ref_349_index_sum_1_req_1); -- 
    -- CP-element group 21 transition  input  output  no-bypass 
    -- predecessors 20 
    -- successors 22 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/final_index_req
      -- 
    partial_sum_1_ca_11033_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_index_sum_1_ack_1, ack => cp_elements(21)); -- 
    final_index_req_11034_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => array_obj_ref_349_offset_inst_req_0); -- 
    -- CP-element group 22 transition  input  output  no-bypass 
    -- predecessors 21 
    -- successors 23 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_base_plus_offset/$entry
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_offset_calculated
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/final_index_ack
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_add_indices/$exit
      -- 
    final_index_ack_11035_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_offset_inst_ack_0, ack => cp_elements(22)); -- 
    sum_rename_req_11039_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => array_obj_ref_349_root_address_inst_req_0); -- 
    -- CP-element group 23 transition  input  no-bypass 
    -- predecessors 22 
    -- successors 10 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_base_plus_offset/$exit
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_root_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_351/array_obj_ref_349_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_11040_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_349_root_address_inst_ack_0, ack => cp_elements(23)); -- 
    -- CP-element group 24 transition  output  bypass 
    -- predecessors 10 
    -- successors 25 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_351/addr_of_350_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_351/addr_of_350_complete/final_reg_req
      -- 
    cp_elements(24) <= cp_elements(10);
    final_reg_req_11044_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => addr_of_350_final_reg_req_0); -- 
    -- CP-element group 25 transition  input  no-bypass 
    -- predecessors 24 
    -- successors 11 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_351/addr_of_350_complete/$exit
      -- 	branch_block_stmt_323/assign_stmt_351/addr_of_350_complete/final_reg_ack
      -- 
    final_reg_ack_11045_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_350_final_reg_ack_0, ack => cp_elements(25)); -- 
    -- CP-element group 26 join  transition  place  bypass 
    -- predecessors 28 11 
    -- successors 29 
    -- members (7) 
      -- 	branch_block_stmt_323/assign_stmt_354/assign_stmt_354_trigger_
      -- 	branch_block_stmt_323/assign_stmt_354/assign_stmt_354_active_
      -- 	branch_block_stmt_323/assign_stmt_354/simple_obj_ref_353_completed_
      -- 	branch_block_stmt_323/assign_stmt_354/$exit
      -- 	branch_block_stmt_323/assign_stmt_354/assign_stmt_354_completed_
      -- 	branch_block_stmt_323/assign_stmt_354__exit__
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370__entry__
      -- 
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(28);
      predecessors(1) <= cp_elements(11);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(26)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 27 transition  output  bypass 
    -- predecessors 11 
    -- successors 28 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_354/simple_obj_ref_353_complete/req
      -- 	branch_block_stmt_323/assign_stmt_354/simple_obj_ref_353_complete/$entry
      -- 
    cp_elements(27) <= cp_elements(11);
    req_11058_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => simple_obj_ref_353_inst_req_0); -- 
    -- CP-element group 28 transition  input  no-bypass 
    -- predecessors 27 
    -- successors 26 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_354/simple_obj_ref_353_complete/ack
      -- 	branch_block_stmt_323/assign_stmt_354/simple_obj_ref_353_complete/$exit
      -- 
    ack_11059_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_353_inst_ack_0, ack => cp_elements(28)); -- 
    -- CP-element group 29 fork  transition  bypass 
    -- predecessors 26 
    -- successors 47 35 31 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/$entry
      -- 
    cp_elements(29) <= cp_elements(26);
    -- CP-element group 30 join  transition  no-bypass 
    -- predecessors 31 34 
    -- successors 58 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_358_completed_
      -- 
    cpelement_group_30 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(31);
      predecessors(1) <= cp_elements(34);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(30)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(30),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 31 fork  transition  bypass 
    -- predecessors 29 
    -- successors 30 32 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_358_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_358_active_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_357_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_357_completed_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_357_active_
      -- 
    cp_elements(31) <= cp_elements(29);
    -- CP-element group 32 join  fork  transition  no-bypass 
    -- predecessors 35 39 31 
    -- successors 40 33 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_trigger_
      -- 
    cpelement_group_32 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(35);
      predecessors(1) <= cp_elements(39);
      predecessors(2) <= cp_elements(31);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(32)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(32),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 33 join  fork  transition  bypass 
    -- predecessors 42 32 
    -- successors 43 34 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_active_
      -- 
    cpelement_group_33 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(42);
      predecessors(1) <= cp_elements(32);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(33)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(33),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 34 join  transition  bypass 
    -- predecessors 44 33 
    -- successors 30 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_completed_
      -- 
    cpelement_group_34 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(44);
      predecessors(1) <= cp_elements(33);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(34)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(34),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 35 fork  transition  bypass 
    -- predecessors 29 
    -- successors 36 32 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_355_completed_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_355_active_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_355_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_address_calculated
      -- 
    cp_elements(35) <= cp_elements(29);
    -- CP-element group 36 transition  output  bypass 
    -- predecessors 35 
    -- successors 37 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_addr_resize/$entry
      -- 
    cp_elements(36) <= cp_elements(35);
    base_resize_req_11082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_356_base_resize_req_0); -- 
    -- CP-element group 37 transition  input  output  no-bypass 
    -- predecessors 36 
    -- successors 38 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_plus_offset/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_address_resized
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_addr_resize/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_11083_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_356_base_resize_ack_0, ack => cp_elements(37)); -- 
    sum_rename_req_11087_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_356_root_address_inst_req_0); -- 
    -- CP-element group 38 transition  input  output  no-bypass 
    -- predecessors 37 
    -- successors 39 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_plus_offset/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_word_addrgen/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_root_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_word_addrgen/root_register_req
      -- 
    sum_rename_ack_11088_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_356_root_address_inst_ack_0, ack => cp_elements(38)); -- 
    root_register_req_11092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => ptr_deref_356_addr_0_req_0); -- 
    -- CP-element group 39 transition  input  no-bypass 
    -- predecessors 38 
    -- successors 32 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_word_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_word_addrgen/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_word_addrgen/root_register_ack
      -- 
    root_register_ack_11093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_356_addr_0_ack_0, ack => cp_elements(39)); -- 
    -- CP-element group 40 transition  output  bypass 
    -- predecessors 32 
    -- successors 41 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/split_req
      -- 
    cp_elements(40) <= cp_elements(32);
    split_req_11097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_356_gather_scatter_req_0); -- 
    -- CP-element group 41 transition  input  output  no-bypass 
    -- predecessors 40 
    -- successors 42 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/word_access/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/split_ack
      -- 
    split_ack_11098_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_356_gather_scatter_ack_0, ack => cp_elements(41)); -- 
    rr_11105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_356_store_0_req_0); -- 
    -- CP-element group 42 transition  input  no-bypass 
    -- predecessors 41 
    -- successors 33 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/word_access/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_request/$exit
      -- 
    ra_11106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_356_store_0_ack_0, ack => cp_elements(42)); -- 
    -- CP-element group 43 transition  output  bypass 
    -- predecessors 33 
    -- successors 44 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/word_access/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/word_access/word_access_0/$entry
      -- 
    cp_elements(43) <= cp_elements(33);
    cr_11116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_356_store_0_req_1); -- 
    -- CP-element group 44 transition  input  no-bypass 
    -- predecessors 43 
    -- successors 34 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/word_access/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/ptr_deref_356_complete/word_access/word_access_0/$exit
      -- 
    ca_11117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_356_store_0_ack_1, ack => cp_elements(44)); -- 
    -- CP-element group 45 join  fork  transition  no-bypass 
    -- predecessors 49 47 
    -- successors 50 46 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_active_
      -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(49);
      predecessors(1) <= cp_elements(47);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(45)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 46 join  fork  transition  bypass 
    -- predecessors 51 45 
    -- successors 52 54 
    -- members (8) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_366_active_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_366_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_364_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_completed_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_366_completed_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_364_active_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_364_completed_
      -- 
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(51);
      predecessors(1) <= cp_elements(45);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(46)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 47 fork  transition  bypass 
    -- predecessors 29 
    -- successors 48 45 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_360_active_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_360_completed_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/simple_obj_ref_360_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_trigger_
      -- 
    cp_elements(47) <= cp_elements(29);
    -- CP-element group 48 transition  output  bypass 
    -- predecessors 47 
    -- successors 49 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Sample/rr
      -- 
    cp_elements(48) <= cp_elements(47);
    rr_11130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => binary_363_inst_req_0); -- 
    -- CP-element group 49 transition  input  no-bypass 
    -- predecessors 48 
    -- successors 45 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Sample/ra
      -- 
    ra_11131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_363_inst_ack_0, ack => cp_elements(49)); -- 
    -- CP-element group 50 transition  output  bypass 
    -- predecessors 45 
    -- successors 51 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Update/cr
      -- 
    cp_elements(50) <= cp_elements(45);
    cr_11135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => binary_363_inst_req_1); -- 
    -- CP-element group 51 transition  input  no-bypass 
    -- predecessors 50 
    -- successors 46 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_363_complete_Update/ca
      -- 
    ca_11136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_363_inst_ack_1, ack => cp_elements(51)); -- 
    -- CP-element group 52 join  fork  transition  bypass 
    -- predecessors 46 55 
    -- successors 56 53 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_active_
      -- 
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(46);
      predecessors(1) <= cp_elements(55);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(52)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 53 join  transition  bypass 
    -- predecessors 57 52 
    -- successors 58 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_370_active_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_completed_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_370_trigger_
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/assign_stmt_370_completed_
      -- 
    cpelement_group_53 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(57);
      predecessors(1) <= cp_elements(52);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(53)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(53),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 54 transition  output  bypass 
    -- predecessors 46 
    -- successors 55 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Sample/rr
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Sample/$entry
      -- 
    cp_elements(54) <= cp_elements(46);
    rr_11149_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => binary_369_inst_req_0); -- 
    -- CP-element group 55 transition  input  no-bypass 
    -- predecessors 54 
    -- successors 52 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Sample/ra
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Sample/$exit
      -- 
    ra_11150_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_369_inst_ack_0, ack => cp_elements(55)); -- 
    -- CP-element group 56 transition  output  bypass 
    -- predecessors 52 
    -- successors 57 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Update/cr
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Update/$entry
      -- 
    cp_elements(56) <= cp_elements(52);
    cr_11154_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => binary_369_inst_req_1); -- 
    -- CP-element group 57 transition  input  no-bypass 
    -- predecessors 56 
    -- successors 53 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Update/ca
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/binary_369_complete_Update/$exit
      -- 
    ca_11155_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_369_inst_ack_1, ack => cp_elements(57)); -- 
    -- CP-element group 58 join  transition  no-bypass 
    -- predecessors 30 53 
    -- successors 1 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_358_to_assign_stmt_370/$exit
      -- 
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(30);
      predecessors(1) <= cp_elements(53);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(58)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 59 transition  bypass 
    -- predecessors 1 
    -- successors 60 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_371_dead_link/$entry
      -- 
    cp_elements(59) <= cp_elements(1);
    -- CP-element group 60 transition  dead  bypass 
    -- predecessors 59 
    -- successors 61 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_371_dead_link/dead_transition
      -- 
    cp_elements(60) <= false;
    -- CP-element group 61 transition  place  bypass 
    -- predecessors 60 
    -- successors 255 
    -- members (4) 
      -- 	branch_block_stmt_323/if_stmt_371_dead_link/$exit
      -- 	branch_block_stmt_323/if_stmt_371__exit__
      -- 	branch_block_stmt_323/merge_stmt_377__entry__
      -- 	branch_block_stmt_323/merge_stmt_377_dead_link/$entry
      -- 
    cp_elements(61) <= cp_elements(60);
    -- CP-element group 62 transition  output  bypass 
    -- predecessors 1 
    -- successors 63 
    -- members (3) 
      -- 	branch_block_stmt_323/if_stmt_371_eval_test/$exit
      -- 	branch_block_stmt_323/if_stmt_371_eval_test/branch_req
      -- 	branch_block_stmt_323/if_stmt_371_eval_test/$entry
      -- 
    cp_elements(62) <= cp_elements(1);
    branch_req_11163_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => if_stmt_371_branch_req_0); -- 
    -- CP-element group 63 branch  place  bypass 
    -- predecessors 62 
    -- successors 64 66 
    -- members (1) 
      -- 	branch_block_stmt_323/simple_obj_ref_372_place
      -- 
    cp_elements(63) <= cp_elements(62);
    -- CP-element group 64 transition  bypass 
    -- predecessors 63 
    -- successors 65 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_371_if_link/$entry
      -- 
    cp_elements(64) <= cp_elements(63);
    -- CP-element group 65 transition  place  input  no-bypass 
    -- predecessors 64 
    -- successors 2 
    -- members (9) 
      -- 	branch_block_stmt_323/if_stmt_371_if_link/if_choice_transition
      -- 	branch_block_stmt_323/if_stmt_371_if_link/$exit
      -- 	branch_block_stmt_323/bb_3_xx_x_crit_edge12x_xi
      -- 	branch_block_stmt_323/merge_stmt_377_PhiAck/dummy
      -- 	branch_block_stmt_323/merge_stmt_377_PhiAck/$exit
      -- 	branch_block_stmt_323/merge_stmt_377_PhiAck/$entry
      -- 	branch_block_stmt_323/bb_3_xx_x_crit_edge12x_xi_PhiReq/$exit
      -- 	branch_block_stmt_323/bb_3_xx_x_crit_edge12x_xi_PhiReq/$entry
      -- 	branch_block_stmt_323/merge_stmt_377_PhiReqMerge
      -- 
    if_choice_transition_11168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_371_branch_ack_1, ack => cp_elements(65)); -- 
    -- CP-element group 66 transition  bypass 
    -- predecessors 63 
    -- successors 67 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_371_else_link/$entry
      -- 
    cp_elements(66) <= cp_elements(63);
    -- CP-element group 67 transition  place  input  output  no-bypass 
    -- predecessors 66 
    -- successors 251 
    -- members (8) 
      -- 	branch_block_stmt_323/bb_3_bb_3
      -- 	branch_block_stmt_323/if_stmt_371_else_link/$exit
      -- 	branch_block_stmt_323/if_stmt_371_else_link/else_choice_transition
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/req
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/$entry
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/$entry
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/$entry
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/$entry
      -- 
    else_choice_transition_11172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_371_branch_ack_0, ack => cp_elements(67)); -- 
    req_11811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => type_cast_344_inst_req_0); -- 
    -- CP-element group 68 join  fork  transition  bypass 
    -- predecessors 71 2 
    -- successors 69 72 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_active_
      -- 
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(71);
      predecessors(1) <= cp_elements(2);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(68)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 69 join  fork  transition  bypass 
    -- predecessors 73 68 
    -- successors 76 74 
    -- members (8) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/assign_stmt_383_active_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/assign_stmt_383_trigger_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/simple_obj_ref_385_active_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/simple_obj_ref_385_trigger_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/simple_obj_ref_385_completed_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_trigger_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/assign_stmt_383_completed_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_completed_
      -- 
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(73);
      predecessors(1) <= cp_elements(68);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(69)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 70 transition  output  bypass 
    -- predecessors 2 
    -- successors 71 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Sample/rr
      -- 
    cp_elements(70) <= cp_elements(2);
    rr_11190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => binary_382_inst_req_0); -- 
    -- CP-element group 71 transition  input  no-bypass 
    -- predecessors 70 
    -- successors 68 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Sample/ra
      -- 
    ra_11191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_382_inst_ack_0, ack => cp_elements(71)); -- 
    -- CP-element group 72 transition  output  bypass 
    -- predecessors 68 
    -- successors 73 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Update/cr
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Update/$entry
      -- 
    cp_elements(72) <= cp_elements(68);
    cr_11195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => binary_382_inst_req_1); -- 
    -- CP-element group 73 transition  input  no-bypass 
    -- predecessors 72 
    -- successors 69 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_382_complete_Update/ca
      -- 
    ca_11196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_382_inst_ack_1, ack => cp_elements(73)); -- 
    -- CP-element group 74 join  fork  transition  no-bypass 
    -- predecessors 77 69 
    -- successors 78 75 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_active_
      -- 
    cpelement_group_74 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(77);
      predecessors(1) <= cp_elements(69);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(74)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(74),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 75 branch  join  transition  place  bypass 
    -- predecessors 79 74 
    -- successors 80 83 
    -- members (7) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/$exit
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_completed_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/assign_stmt_389_active_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/assign_stmt_389_trigger_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/assign_stmt_389_completed_
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389__exit__
      -- 	branch_block_stmt_323/if_stmt_390__entry__
      -- 
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(79);
      predecessors(1) <= cp_elements(74);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(75)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 76 transition  output  bypass 
    -- predecessors 69 
    -- successors 77 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Sample/rr
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Sample/$entry
      -- 
    cp_elements(76) <= cp_elements(69);
    rr_11209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => binary_388_inst_req_0); -- 
    -- CP-element group 77 transition  input  no-bypass 
    -- predecessors 76 
    -- successors 74 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Sample/ra
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Sample/$exit
      -- 
    ra_11210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_388_inst_ack_0, ack => cp_elements(77)); -- 
    -- CP-element group 78 transition  output  bypass 
    -- predecessors 74 
    -- successors 79 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Update/cr
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Update/$entry
      -- 
    cp_elements(78) <= cp_elements(74);
    cr_11214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => binary_388_inst_req_1); -- 
    -- CP-element group 79 transition  input  no-bypass 
    -- predecessors 78 
    -- successors 75 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_383_to_assign_stmt_389/binary_388_complete_Update/ca
      -- 
    ca_11215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_388_inst_ack_1, ack => cp_elements(79)); -- 
    -- CP-element group 80 transition  bypass 
    -- predecessors 75 
    -- successors 81 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_390_dead_link/$entry
      -- 
    cp_elements(80) <= cp_elements(75);
    -- CP-element group 81 transition  dead  bypass 
    -- predecessors 80 
    -- successors 82 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_390_dead_link/dead_transition
      -- 
    cp_elements(81) <= false;
    -- CP-element group 82 transition  place  bypass 
    -- predecessors 81 
    -- successors 257 
    -- members (4) 
      -- 	branch_block_stmt_323/if_stmt_390_dead_link/$exit
      -- 	branch_block_stmt_323/if_stmt_390__exit__
      -- 	branch_block_stmt_323/merge_stmt_396__entry__
      -- 	branch_block_stmt_323/merge_stmt_396_dead_link/$entry
      -- 
    cp_elements(82) <= cp_elements(81);
    -- CP-element group 83 transition  output  bypass 
    -- predecessors 75 
    -- successors 84 
    -- members (3) 
      -- 	branch_block_stmt_323/if_stmt_390_eval_test/$entry
      -- 	branch_block_stmt_323/if_stmt_390_eval_test/branch_req
      -- 	branch_block_stmt_323/if_stmt_390_eval_test/$exit
      -- 
    cp_elements(83) <= cp_elements(75);
    branch_req_11223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => if_stmt_390_branch_req_0); -- 
    -- CP-element group 84 branch  place  bypass 
    -- predecessors 83 
    -- successors 85 87 
    -- members (1) 
      -- 	branch_block_stmt_323/simple_obj_ref_391_place
      -- 
    cp_elements(84) <= cp_elements(83);
    -- CP-element group 85 transition  bypass 
    -- predecessors 84 
    -- successors 86 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_390_if_link/$entry
      -- 
    cp_elements(85) <= cp_elements(84);
    -- CP-element group 86 transition  place  input  output  no-bypass 
    -- predecessors 85 
    -- successors 264 
    -- members (22) 
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnphx_xix_xpreheader
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_req
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/ack
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/req
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/$exit
      -- 	branch_block_stmt_323/if_stmt_390_if_link/$exit
      -- 	branch_block_stmt_323/if_stmt_390_if_link/if_choice_transition
      -- 	branch_block_stmt_323/merge_stmt_406__exit__
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/phi_stmt_409/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xix_xpreheader_bbx_xnphx_xi_PhiReq/$entry
      -- 	branch_block_stmt_323/merge_stmt_406_PhiAck/dummy
      -- 	branch_block_stmt_323/merge_stmt_406_PhiAck/$exit
      -- 	branch_block_stmt_323/merge_stmt_406_PhiAck/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnphx_xix_xpreheader_PhiReq/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnphx_xix_xpreheader_PhiReq/$entry
      -- 	branch_block_stmt_323/merge_stmt_406_PhiReqMerge
      -- 
    if_choice_transition_11228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_390_branch_ack_1, ack => cp_elements(86)); -- 
    phi_stmt_409_req_11907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => phi_stmt_409_req_1); -- 
    -- CP-element group 87 transition  bypass 
    -- predecessors 84 
    -- successors 88 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_390_else_link/$entry
      -- 
    cp_elements(87) <= cp_elements(84);
    -- CP-element group 88 transition  place  input  output  no-bypass 
    -- predecessors 87 
    -- successors 259 
    -- members (8) 
      -- 	branch_block_stmt_323/if_stmt_390_else_link/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge
      -- 	branch_block_stmt_323/if_stmt_390_else_link/else_choice_transition
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/req
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/$entry
      -- 
    else_choice_transition_11232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_390_branch_ack_0, ack => cp_elements(88)); -- 
    req_11877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => type_cast_400_inst_req_0); -- 
    -- CP-element group 89 fork  transition  bypass 
    -- predecessors 270 
    -- successors 90 94 98 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_432/$entry
      -- 
    cp_elements(89) <= cp_elements(270);
    -- CP-element group 90 transition  bypass 
    -- predecessors 89 
    -- successors 91 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_432/addr_of_431_trigger_
      -- 
    cp_elements(90) <= cp_elements(89);
    -- CP-element group 91 join  fork  transition  bypass 
    -- predecessors 90 104 
    -- successors 92 105 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_432/addr_of_431_active_
      -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(90);
      predecessors(1) <= cp_elements(104);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(91)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 92 join  fork  transition  place  no-bypass 
    -- predecessors 91 106 
    -- successors 107 108 
    -- members (10) 
      -- 	branch_block_stmt_323/assign_stmt_432/addr_of_431_completed_
      -- 	branch_block_stmt_323/assign_stmt_435/$entry
      -- 	branch_block_stmt_323/assign_stmt_435/simple_obj_ref_434_active_
      -- 	branch_block_stmt_323/assign_stmt_432/assign_stmt_432_trigger_
      -- 	branch_block_stmt_323/assign_stmt_432/assign_stmt_432_completed_
      -- 	branch_block_stmt_323/assign_stmt_432/assign_stmt_432_active_
      -- 	branch_block_stmt_323/assign_stmt_435/simple_obj_ref_434_trigger_
      -- 	branch_block_stmt_323/assign_stmt_432/$exit
      -- 	branch_block_stmt_323/assign_stmt_432__exit__
      -- 	branch_block_stmt_323/assign_stmt_435__entry__
      -- 
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(91);
      predecessors(1) <= cp_elements(106);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(92)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 93 join  transition  output  bypass 
    -- predecessors 97 100 
    -- successors 101 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_indices_scaled
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/$entry
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(97);
      predecessors(1) <= cp_elements(100);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(93)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_11282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => array_obj_ref_430_index_sum_1_req_0); -- 
    -- CP-element group 94 transition  output  bypass 
    -- predecessors 89 
    -- successors 95 
    -- members (6) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_0/index_resize_req
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_432/simple_obj_ref_428_completed_
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_computed_0
      -- 	branch_block_stmt_323/assign_stmt_432/simple_obj_ref_428_active_
      -- 	branch_block_stmt_323/assign_stmt_432/simple_obj_ref_428_trigger_
      -- 
    cp_elements(94) <= cp_elements(89);
    index_resize_req_11255_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => array_obj_ref_430_index_0_resize_req_0); -- 
    -- CP-element group 95 transition  input  output  no-bypass 
    -- predecessors 94 
    -- successors 96 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resized_0
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_0/scale_rr
      -- 
    index_resize_ack_11256_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_0_resize_ack_0, ack => cp_elements(95)); -- 
    scale_rr_11260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => array_obj_ref_430_index_0_scale_req_0); -- 
    -- CP-element group 96 transition  input  output  no-bypass 
    -- predecessors 95 
    -- successors 97 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_0/scale_ra
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_0/scale_cr
      -- 
    scale_ra_11261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_0_scale_ack_0, ack => cp_elements(96)); -- 
    scale_cr_11262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => array_obj_ref_430_index_0_scale_req_1); -- 
    -- CP-element group 97 transition  input  no-bypass 
    -- predecessors 96 
    -- successors 93 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_0/scale_ca
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_0/$exit
      -- 
    scale_ca_11263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_0_scale_ack_1, ack => cp_elements(97)); -- 
    -- CP-element group 98 transition  output  bypass 
    -- predecessors 89 
    -- successors 99 
    -- members (6) 
      -- 	branch_block_stmt_323/assign_stmt_432/simple_obj_ref_429_completed_
      -- 	branch_block_stmt_323/assign_stmt_432/simple_obj_ref_429_active_
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_1/$entry
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_computed_1
      -- 	branch_block_stmt_323/assign_stmt_432/simple_obj_ref_429_trigger_
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_1/index_resize_req
      -- 
    cp_elements(98) <= cp_elements(89);
    index_resize_req_11272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => array_obj_ref_430_index_1_resize_req_0); -- 
    -- CP-element group 99 transition  input  output  no-bypass 
    -- predecessors 98 
    -- successors 100 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_1/$exit
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_resized_1
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_1/$entry
      -- 
    index_resize_ack_11273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_1_resize_ack_0, ack => cp_elements(99)); -- 
    scale_rename_req_11277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => array_obj_ref_430_index_1_rename_req_0); -- 
    -- CP-element group 100 transition  input  no-bypass 
    -- predecessors 99 
    -- successors 93 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_index_scale_1/$exit
      -- 
    scale_rename_ack_11278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_1_rename_ack_0, ack => cp_elements(100)); -- 
    -- CP-element group 101 transition  input  output  no-bypass 
    -- predecessors 93 
    -- successors 102 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_11283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_sum_1_ack_0, ack => cp_elements(101)); -- 
    partial_sum_1_cr_11284_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => array_obj_ref_430_index_sum_1_req_1); -- 
    -- CP-element group 102 transition  input  output  no-bypass 
    -- predecessors 101 
    -- successors 103 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/final_index_req
      -- 
    partial_sum_1_ca_11285_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_sum_1_ack_1, ack => cp_elements(102)); -- 
    final_index_req_11286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => array_obj_ref_430_offset_inst_req_0); -- 
    -- CP-element group 103 transition  input  output  no-bypass 
    -- predecessors 102 
    -- successors 104 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/final_index_ack
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_offset_calculated
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_base_plus_offset/$entry
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_add_indices/$exit
      -- 
    final_index_ack_11287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_offset_inst_ack_0, ack => cp_elements(103)); -- 
    sum_rename_req_11291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => array_obj_ref_430_root_address_inst_req_0); -- 
    -- CP-element group 104 transition  input  no-bypass 
    -- predecessors 103 
    -- successors 91 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_root_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_base_plus_offset/$exit
      -- 	branch_block_stmt_323/assign_stmt_432/array_obj_ref_430_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_11292_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_root_address_inst_ack_0, ack => cp_elements(104)); -- 
    -- CP-element group 105 transition  output  bypass 
    -- predecessors 91 
    -- successors 106 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_432/addr_of_431_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_432/addr_of_431_complete/final_reg_req
      -- 
    cp_elements(105) <= cp_elements(91);
    final_reg_req_11296_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => addr_of_431_final_reg_req_0); -- 
    -- CP-element group 106 transition  input  no-bypass 
    -- predecessors 105 
    -- successors 92 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_432/addr_of_431_complete/final_reg_ack
      -- 	branch_block_stmt_323/assign_stmt_432/addr_of_431_complete/$exit
      -- 
    final_reg_ack_11297_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_431_final_reg_ack_0, ack => cp_elements(106)); -- 
    -- CP-element group 107 join  transition  place  bypass 
    -- predecessors 92 109 
    -- successors 110 
    -- members (7) 
      -- 	branch_block_stmt_323/assign_stmt_435/assign_stmt_435_completed_
      -- 	branch_block_stmt_323/assign_stmt_435/$exit
      -- 	branch_block_stmt_323/assign_stmt_435/assign_stmt_435_trigger_
      -- 	branch_block_stmt_323/assign_stmt_435/assign_stmt_435_active_
      -- 	branch_block_stmt_323/assign_stmt_435/simple_obj_ref_434_completed_
      -- 	branch_block_stmt_323/assign_stmt_435__exit__
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451__entry__
      -- 
    cpelement_group_107 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(92);
      predecessors(1) <= cp_elements(109);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(107)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(107),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 108 transition  output  bypass 
    -- predecessors 92 
    -- successors 109 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_435/simple_obj_ref_434_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_435/simple_obj_ref_434_complete/req
      -- 
    cp_elements(108) <= cp_elements(92);
    req_11310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => simple_obj_ref_434_inst_req_0); -- 
    -- CP-element group 109 transition  input  no-bypass 
    -- predecessors 108 
    -- successors 107 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_435/simple_obj_ref_434_complete/ack
      -- 	branch_block_stmt_323/assign_stmt_435/simple_obj_ref_434_complete/$exit
      -- 
    ack_11311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_434_inst_ack_0, ack => cp_elements(109)); -- 
    -- CP-element group 110 fork  transition  bypass 
    -- predecessors 107 
    -- successors 112 116 128 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/$entry
      -- 
    cp_elements(110) <= cp_elements(107);
    -- CP-element group 111 join  transition  no-bypass 
    -- predecessors 112 115 
    -- successors 139 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_439_completed_
      -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(112);
      predecessors(1) <= cp_elements(115);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(111)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 112 fork  transition  bypass 
    -- predecessors 110 
    -- successors 111 113 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_439_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_439_active_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_438_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_438_active_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_438_completed_
      -- 
    cp_elements(112) <= cp_elements(110);
    -- CP-element group 113 join  fork  transition  no-bypass 
    -- predecessors 112 116 120 
    -- successors 114 121 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_trigger_
      -- 
    cpelement_group_113 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(112);
      predecessors(1) <= cp_elements(116);
      predecessors(2) <= cp_elements(120);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(113)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 114 join  fork  transition  bypass 
    -- predecessors 113 123 
    -- successors 115 124 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_active_
      -- 
    cpelement_group_114 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(113);
      predecessors(1) <= cp_elements(123);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(114)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(114),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 115 join  transition  bypass 
    -- predecessors 114 125 
    -- successors 111 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_completed_
      -- 
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(114);
      predecessors(1) <= cp_elements(125);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(115)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 116 fork  transition  bypass 
    -- predecessors 110 
    -- successors 113 117 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_436_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_436_active_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_436_completed_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_address_calculated
      -- 
    cp_elements(116) <= cp_elements(110);
    -- CP-element group 117 transition  output  bypass 
    -- predecessors 116 
    -- successors 118 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_addr_resize/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_addr_resize/base_resize_req
      -- 
    cp_elements(117) <= cp_elements(116);
    base_resize_req_11334_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_437_base_resize_req_0); -- 
    -- CP-element group 118 transition  input  output  no-bypass 
    -- predecessors 117 
    -- successors 119 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_address_resized
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_plus_offset/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_addr_resize/$exit
      -- 
    base_resize_ack_11335_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_437_base_resize_ack_0, ack => cp_elements(118)); -- 
    sum_rename_req_11339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => ptr_deref_437_root_address_inst_req_0); -- 
    -- CP-element group 119 transition  input  output  no-bypass 
    -- predecessors 118 
    -- successors 120 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_word_addrgen/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_word_addrgen/root_register_req
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_root_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_base_plus_offset/$exit
      -- 
    sum_rename_ack_11340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_437_root_address_inst_ack_0, ack => cp_elements(119)); -- 
    root_register_req_11344_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => ptr_deref_437_addr_0_req_0); -- 
    -- CP-element group 120 transition  input  no-bypass 
    -- predecessors 119 
    -- successors 113 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_word_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_word_addrgen/root_register_ack
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_word_addrgen/$exit
      -- 
    root_register_ack_11345_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_437_addr_0_ack_0, ack => cp_elements(120)); -- 
    -- CP-element group 121 transition  output  bypass 
    -- predecessors 113 
    -- successors 122 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/split_req
      -- 
    cp_elements(121) <= cp_elements(113);
    split_req_11349_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => ptr_deref_437_gather_scatter_req_0); -- 
    -- CP-element group 122 transition  input  output  no-bypass 
    -- predecessors 121 
    -- successors 123 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/split_ack
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/word_access/$entry
      -- 
    split_ack_11350_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_437_gather_scatter_ack_0, ack => cp_elements(122)); -- 
    rr_11357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_437_store_0_req_0); -- 
    -- CP-element group 123 transition  input  no-bypass 
    -- predecessors 122 
    -- successors 114 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/$exit
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_request/word_access/$exit
      -- 
    ra_11358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_437_store_0_ack_0, ack => cp_elements(123)); -- 
    -- CP-element group 124 transition  output  bypass 
    -- predecessors 114 
    -- successors 125 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/word_access/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/word_access/word_access_0/$entry
      -- 
    cp_elements(124) <= cp_elements(114);
    cr_11368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => ptr_deref_437_store_0_req_1); -- 
    -- CP-element group 125 transition  input  no-bypass 
    -- predecessors 124 
    -- successors 115 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/$exit
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/ptr_deref_437_complete/word_access/$exit
      -- 
    ca_11369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_437_store_0_ack_1, ack => cp_elements(125)); -- 
    -- CP-element group 126 join  fork  transition  no-bypass 
    -- predecessors 128 130 
    -- successors 127 131 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_active_
      -- 
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(128);
      predecessors(1) <= cp_elements(130);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(126)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 127 join  fork  transition  bypass 
    -- predecessors 126 132 
    -- successors 133 135 
    -- members (8) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_445_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_445_active_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_445_completed_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_447_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_447_active_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_completed_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_447_completed_
      -- 
    cpelement_group_127 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(126);
      predecessors(1) <= cp_elements(132);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(127)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(127),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 128 fork  transition  bypass 
    -- predecessors 110 
    -- successors 126 129 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_441_active_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_441_completed_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/simple_obj_ref_441_trigger_
      -- 
    cp_elements(128) <= cp_elements(110);
    -- CP-element group 129 transition  output  bypass 
    -- predecessors 128 
    -- successors 130 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Sample/rr
      -- 
    cp_elements(129) <= cp_elements(128);
    rr_11382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => binary_444_inst_req_0); -- 
    -- CP-element group 130 transition  input  no-bypass 
    -- predecessors 129 
    -- successors 126 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Sample/ra
      -- 
    ra_11383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_444_inst_ack_0, ack => cp_elements(130)); -- 
    -- CP-element group 131 transition  output  bypass 
    -- predecessors 126 
    -- successors 132 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Update/cr
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Update/$entry
      -- 
    cp_elements(131) <= cp_elements(126);
    cr_11387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => binary_444_inst_req_1); -- 
    -- CP-element group 132 transition  input  no-bypass 
    -- predecessors 131 
    -- successors 127 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Update/ca
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_444_complete_Update/$exit
      -- 
    ca_11388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_444_inst_ack_1, ack => cp_elements(132)); -- 
    -- CP-element group 133 join  fork  transition  bypass 
    -- predecessors 127 136 
    -- successors 134 137 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_active_
      -- 
    cpelement_group_133 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(127);
      predecessors(1) <= cp_elements(136);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(133)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(133),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 134 join  transition  no-bypass 
    -- predecessors 133 138 
    -- successors 139 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_451_trigger_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_451_completed_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_completed_
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/assign_stmt_451_active_
      -- 
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(133);
      predecessors(1) <= cp_elements(138);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(134)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 135 transition  output  bypass 
    -- predecessors 127 
    -- successors 136 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Sample/rr
      -- 
    cp_elements(135) <= cp_elements(127);
    rr_11401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => binary_450_inst_req_0); -- 
    -- CP-element group 136 transition  input  no-bypass 
    -- predecessors 135 
    -- successors 133 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Sample/ra
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Sample/$exit
      -- 
    ra_11402_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_450_inst_ack_0, ack => cp_elements(136)); -- 
    -- CP-element group 137 transition  output  bypass 
    -- predecessors 133 
    -- successors 138 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Update/cr
      -- 
    cp_elements(137) <= cp_elements(133);
    cr_11406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(137), ack => binary_450_inst_req_1); -- 
    -- CP-element group 138 transition  input  no-bypass 
    -- predecessors 137 
    -- successors 134 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/binary_450_complete_Update/ca
      -- 
    ca_11407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_450_inst_ack_1, ack => cp_elements(138)); -- 
    -- CP-element group 139 join  transition  no-bypass 
    -- predecessors 111 134 
    -- successors 4 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_439_to_assign_stmt_451/$exit
      -- 
    cpelement_group_139 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(111);
      predecessors(1) <= cp_elements(134);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(139)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(139),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 140 transition  bypass 
    -- predecessors 4 
    -- successors 141 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_452_dead_link/$entry
      -- 
    cp_elements(140) <= cp_elements(4);
    -- CP-element group 141 transition  dead  bypass 
    -- predecessors 140 
    -- successors 142 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_452_dead_link/dead_transition
      -- 
    cp_elements(141) <= false;
    -- CP-element group 142 transition  place  bypass 
    -- predecessors 141 
    -- successors 271 
    -- members (4) 
      -- 	branch_block_stmt_323/merge_stmt_458_dead_link/$entry
      -- 	branch_block_stmt_323/if_stmt_452_dead_link/$exit
      -- 	branch_block_stmt_323/if_stmt_452__exit__
      -- 	branch_block_stmt_323/merge_stmt_458__entry__
      -- 
    cp_elements(142) <= cp_elements(141);
    -- CP-element group 143 transition  output  bypass 
    -- predecessors 4 
    -- successors 144 
    -- members (3) 
      -- 	branch_block_stmt_323/if_stmt_452_eval_test/branch_req
      -- 	branch_block_stmt_323/if_stmt_452_eval_test/$entry
      -- 	branch_block_stmt_323/if_stmt_452_eval_test/$exit
      -- 
    cp_elements(143) <= cp_elements(4);
    branch_req_11415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(143), ack => if_stmt_452_branch_req_0); -- 
    -- CP-element group 144 branch  place  bypass 
    -- predecessors 143 
    -- successors 145 147 
    -- members (1) 
      -- 	branch_block_stmt_323/simple_obj_ref_453_place
      -- 
    cp_elements(144) <= cp_elements(143);
    -- CP-element group 145 transition  bypass 
    -- predecessors 144 
    -- successors 146 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_452_if_link/$entry
      -- 
    cp_elements(145) <= cp_elements(144);
    -- CP-element group 146 transition  place  input  no-bypass 
    -- predecessors 145 
    -- successors 5 
    -- members (9) 
      -- 	branch_block_stmt_323/bb_8_xx_x_crit_edgex_xi
      -- 	branch_block_stmt_323/bb_8_xx_x_crit_edgex_xi_PhiReq/$entry
      -- 	branch_block_stmt_323/if_stmt_452_if_link/$exit
      -- 	branch_block_stmt_323/if_stmt_452_if_link/if_choice_transition
      -- 	branch_block_stmt_323/merge_stmt_458_PhiAck/dummy
      -- 	branch_block_stmt_323/merge_stmt_458_PhiAck/$exit
      -- 	branch_block_stmt_323/merge_stmt_458_PhiReqMerge
      -- 	branch_block_stmt_323/merge_stmt_458_PhiAck/$entry
      -- 	branch_block_stmt_323/bb_8_xx_x_crit_edgex_xi_PhiReq/$exit
      -- 
    if_choice_transition_11420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_452_branch_ack_1, ack => cp_elements(146)); -- 
    -- CP-element group 147 transition  bypass 
    -- predecessors 144 
    -- successors 148 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_452_else_link/$entry
      -- 
    cp_elements(147) <= cp_elements(144);
    -- CP-element group 148 transition  place  input  output  no-bypass 
    -- predecessors 147 
    -- successors 267 
    -- members (8) 
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/$entry
      -- 	branch_block_stmt_323/bb_8_bb_8
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/$entry
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/$entry
      -- 	branch_block_stmt_323/if_stmt_452_else_link/$exit
      -- 	branch_block_stmt_323/if_stmt_452_else_link/else_choice_transition
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/$entry
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/req
      -- 
    else_choice_transition_11424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_452_branch_ack_0, ack => cp_elements(148)); -- 
    req_11940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => type_cast_425_inst_req_0); -- 
    -- CP-element group 149 join  fork  transition  bypass 
    -- predecessors 152 5 
    -- successors 150 153 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_active_
      -- 
    cpelement_group_149 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(152);
      predecessors(1) <= cp_elements(5);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(149)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(149),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 150 join  fork  transition  bypass 
    -- predecessors 149 154 
    -- successors 155 157 
    -- members (8) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_trigger_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/simple_obj_ref_466_trigger_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/simple_obj_ref_466_active_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/simple_obj_ref_466_completed_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_completed_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/assign_stmt_464_trigger_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/assign_stmt_464_active_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/assign_stmt_464_completed_
      -- 
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(149);
      predecessors(1) <= cp_elements(154);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(150)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 151 transition  output  bypass 
    -- predecessors 5 
    -- successors 152 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Sample/rr
      -- 
    cp_elements(151) <= cp_elements(5);
    rr_11442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => binary_463_inst_req_0); -- 
    -- CP-element group 152 transition  input  no-bypass 
    -- predecessors 151 
    -- successors 149 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Sample/ra
      -- 
    ra_11443_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_463_inst_ack_0, ack => cp_elements(152)); -- 
    -- CP-element group 153 transition  output  bypass 
    -- predecessors 149 
    -- successors 154 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Update/cr
      -- 
    cp_elements(153) <= cp_elements(149);
    cr_11447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => binary_463_inst_req_1); -- 
    -- CP-element group 154 transition  input  no-bypass 
    -- predecessors 153 
    -- successors 150 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_463_complete_Update/ca
      -- 
    ca_11448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_463_inst_ack_1, ack => cp_elements(154)); -- 
    -- CP-element group 155 join  fork  transition  no-bypass 
    -- predecessors 150 158 
    -- successors 156 159 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_active_
      -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(150);
      predecessors(1) <= cp_elements(158);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(155)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 156 branch  join  transition  place  no-bypass 
    -- predecessors 155 160 
    -- successors 161 164 
    -- members (7) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/assign_stmt_470_trigger_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/assign_stmt_470_active_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/assign_stmt_470_completed_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_completed_
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/$exit
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470__exit__
      -- 	branch_block_stmt_323/if_stmt_471__entry__
      -- 
    cpelement_group_156 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(155);
      predecessors(1) <= cp_elements(160);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(156)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(156),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 157 transition  output  bypass 
    -- predecessors 150 
    -- successors 158 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Sample/rr
      -- 
    cp_elements(157) <= cp_elements(150);
    rr_11461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => binary_469_inst_req_0); -- 
    -- CP-element group 158 transition  input  no-bypass 
    -- predecessors 157 
    -- successors 155 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Sample/ra
      -- 
    ra_11462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_469_inst_ack_0, ack => cp_elements(158)); -- 
    -- CP-element group 159 transition  output  bypass 
    -- predecessors 155 
    -- successors 160 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Update/cr
      -- 
    cp_elements(159) <= cp_elements(155);
    cr_11466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(159), ack => binary_469_inst_req_1); -- 
    -- CP-element group 160 transition  input  no-bypass 
    -- predecessors 159 
    -- successors 156 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_464_to_assign_stmt_470/binary_469_complete_Update/ca
      -- 
    ca_11467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_469_inst_ack_1, ack => cp_elements(160)); -- 
    -- CP-element group 161 transition  bypass 
    -- predecessors 156 
    -- successors 162 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_471_dead_link/$entry
      -- 
    cp_elements(161) <= cp_elements(156);
    -- CP-element group 162 transition  dead  bypass 
    -- predecessors 161 
    -- successors 163 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_471_dead_link/dead_transition
      -- 
    cp_elements(162) <= false;
    -- CP-element group 163 transition  place  bypass 
    -- predecessors 162 
    -- successors 273 
    -- members (4) 
      -- 	branch_block_stmt_323/if_stmt_471__exit__
      -- 	branch_block_stmt_323/merge_stmt_477__entry__
      -- 	branch_block_stmt_323/if_stmt_471_dead_link/$exit
      -- 	branch_block_stmt_323/merge_stmt_477_dead_link/$entry
      -- 
    cp_elements(163) <= cp_elements(162);
    -- CP-element group 164 transition  output  bypass 
    -- predecessors 156 
    -- successors 165 
    -- members (3) 
      -- 	branch_block_stmt_323/if_stmt_471_eval_test/$entry
      -- 	branch_block_stmt_323/if_stmt_471_eval_test/$exit
      -- 	branch_block_stmt_323/if_stmt_471_eval_test/branch_req
      -- 
    cp_elements(164) <= cp_elements(156);
    branch_req_11475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => if_stmt_471_branch_req_0); -- 
    -- CP-element group 165 branch  place  bypass 
    -- predecessors 164 
    -- successors 166 168 
    -- members (1) 
      -- 	branch_block_stmt_323/simple_obj_ref_472_place
      -- 
    cp_elements(165) <= cp_elements(164);
    -- CP-element group 166 transition  bypass 
    -- predecessors 165 
    -- successors 167 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_471_if_link/$entry
      -- 
    cp_elements(166) <= cp_elements(165);
    -- CP-element group 167 transition  place  input  no-bypass 
    -- predecessors 166 
    -- successors 6 
    -- members (9) 
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_get_inputx_xexit
      -- 	branch_block_stmt_323/merge_stmt_477_PhiAck/$entry
      -- 	branch_block_stmt_323/merge_stmt_477_PhiAck/dummy
      -- 	branch_block_stmt_323/merge_stmt_477_PhiAck/$exit
      -- 	branch_block_stmt_323/if_stmt_471_if_link/$exit
      -- 	branch_block_stmt_323/if_stmt_471_if_link/if_choice_transition
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_get_inputx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_get_inputx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_323/merge_stmt_477_PhiReqMerge
      -- 
    if_choice_transition_11480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_471_branch_ack_1, ack => cp_elements(167)); -- 
    -- CP-element group 168 transition  bypass 
    -- predecessors 165 
    -- successors 169 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_471_else_link/$entry
      -- 
    cp_elements(168) <= cp_elements(165);
    -- CP-element group 169 transition  place  input  output  no-bypass 
    -- predecessors 168 
    -- successors 263 
    -- members (8) 
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/req
      -- 	branch_block_stmt_323/if_stmt_471_else_link/$exit
      -- 	branch_block_stmt_323/if_stmt_471_else_link/else_choice_transition
      -- 
    else_choice_transition_11484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_471_branch_ack_0, ack => cp_elements(169)); -- 
    req_11920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(169), ack => type_cast_412_inst_req_0); -- 
    -- CP-element group 170 transition  input  output  no-bypass 
    -- predecessors 6 
    -- successors 171 
    -- members (5) 
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_active_
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_start/$exit
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_start/cra
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_complete/$entry
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_complete/ccr
      -- 
    cra_11498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_478_call_ack_0, ack => cp_elements(170)); -- 
    ccr_11502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => call_stmt_478_call_req_1); -- 
    -- CP-element group 171 transition  place  input  output  no-bypass 
    -- predecessors 170 
    -- successors 276 
    -- members (18) 
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/$exit
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/$exit
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/$entry
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/$entry
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1
      -- 	branch_block_stmt_323/call_stmt_478__exit__
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/ack
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/$entry
      -- 	branch_block_stmt_323/call_stmt_478/$exit
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_call_complete
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_completed_
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_complete/$exit
      -- 	branch_block_stmt_323/call_stmt_478/call_stmt_478_complete/cca
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/$exit
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/req
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/$exit
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_req
      -- 	branch_block_stmt_323/get_inputx_xexit_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/$entry
      -- 
    cca_11503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_478_call_ack_1, ack => cp_elements(171)); -- 
    phi_stmt_481_req_12001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => phi_stmt_481_req_0); -- 
    -- CP-element group 172 fork  transition  bypass 
    -- predecessors 282 
    -- successors 173 177 181 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/$entry
      -- 
    cp_elements(172) <= cp_elements(282);
    -- CP-element group 173 transition  bypass 
    -- predecessors 172 
    -- successors 174 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/addr_of_503_trigger_
      -- 
    cp_elements(173) <= cp_elements(172);
    -- CP-element group 174 join  fork  transition  bypass 
    -- predecessors 173 187 
    -- successors 175 188 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/addr_of_503_active_
      -- 
    cpelement_group_174 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(173);
      predecessors(1) <= cp_elements(187);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(174)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(174),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 175 join  transition  output  no-bypass 
    -- predecessors 174 189 
    -- successors 192 
    -- members (10) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/assign_stmt_504_trigger_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/assign_stmt_504_active_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/assign_stmt_504_completed_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/addr_of_503_completed_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_506_trigger_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_506_active_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_506_completed_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_addr_resize/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_addr_resize/base_resize_req
      -- 
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(174);
      predecessors(1) <= cp_elements(189);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(175)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_11583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(175), ack => ptr_deref_507_base_resize_req_0); -- 
    -- CP-element group 176 join  transition  output  bypass 
    -- predecessors 180 183 
    -- successors 184 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_indices_scaled
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(180);
      predecessors(1) <= cp_elements(183);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(176)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_11551_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => array_obj_ref_502_index_sum_1_req_0); -- 
    -- CP-element group 177 transition  output  bypass 
    -- predecessors 172 
    -- successors 178 
    -- members (6) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_computed_0
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_500_trigger_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_500_active_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_500_completed_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_0/index_resize_req
      -- 
    cp_elements(177) <= cp_elements(172);
    index_resize_req_11524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => array_obj_ref_502_index_0_resize_req_0); -- 
    -- CP-element group 178 transition  input  output  no-bypass 
    -- predecessors 177 
    -- successors 179 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resized_0
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_0/scale_rr
      -- 
    index_resize_ack_11525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_index_0_resize_ack_0, ack => cp_elements(178)); -- 
    scale_rr_11529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => array_obj_ref_502_index_0_scale_req_0); -- 
    -- CP-element group 179 transition  input  output  no-bypass 
    -- predecessors 178 
    -- successors 180 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_0/scale_ra
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_0/scale_cr
      -- 
    scale_ra_11530_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_index_0_scale_ack_0, ack => cp_elements(179)); -- 
    scale_cr_11531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => array_obj_ref_502_index_0_scale_req_1); -- 
    -- CP-element group 180 transition  input  no-bypass 
    -- predecessors 179 
    -- successors 176 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_0/scale_ca
      -- 
    scale_ca_11532_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_index_0_scale_ack_1, ack => cp_elements(180)); -- 
    -- CP-element group 181 transition  output  bypass 
    -- predecessors 172 
    -- successors 182 
    -- members (6) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_computed_1
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_501_trigger_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_501_active_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/simple_obj_ref_501_completed_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_1/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_1/index_resize_req
      -- 
    cp_elements(181) <= cp_elements(172);
    index_resize_req_11541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => array_obj_ref_502_index_1_resize_req_0); -- 
    -- CP-element group 182 transition  input  output  no-bypass 
    -- predecessors 181 
    -- successors 183 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resized_1
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_1/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_1/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_11542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_index_1_resize_ack_0, ack => cp_elements(182)); -- 
    scale_rename_req_11546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(182), ack => array_obj_ref_502_index_1_rename_req_0); -- 
    -- CP-element group 183 transition  input  no-bypass 
    -- predecessors 182 
    -- successors 176 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_1/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_11547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_index_1_rename_ack_0, ack => cp_elements(183)); -- 
    -- CP-element group 184 transition  input  output  no-bypass 
    -- predecessors 176 
    -- successors 185 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_11552_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_index_sum_1_ack_0, ack => cp_elements(184)); -- 
    partial_sum_1_cr_11553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(184), ack => array_obj_ref_502_index_sum_1_req_1); -- 
    -- CP-element group 185 transition  input  output  no-bypass 
    -- predecessors 184 
    -- successors 186 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/final_index_req
      -- 
    partial_sum_1_ca_11554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_index_sum_1_ack_1, ack => cp_elements(185)); -- 
    final_index_req_11555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => array_obj_ref_502_offset_inst_req_0); -- 
    -- CP-element group 186 transition  input  output  no-bypass 
    -- predecessors 185 
    -- successors 187 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_offset_calculated
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_add_indices/final_index_ack
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_base_plus_offset/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_11556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_offset_inst_ack_0, ack => cp_elements(186)); -- 
    sum_rename_req_11560_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => array_obj_ref_502_root_address_inst_req_0); -- 
    -- CP-element group 187 transition  input  no-bypass 
    -- predecessors 186 
    -- successors 174 
    -- members (3) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_root_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_base_plus_offset/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/array_obj_ref_502_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_11561_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_502_root_address_inst_ack_0, ack => cp_elements(187)); -- 
    -- CP-element group 188 transition  output  bypass 
    -- predecessors 174 
    -- successors 189 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/addr_of_503_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/addr_of_503_complete/final_reg_req
      -- 
    cp_elements(188) <= cp_elements(174);
    final_reg_req_11565_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => addr_of_503_final_reg_req_0); -- 
    -- CP-element group 189 transition  input  no-bypass 
    -- predecessors 188 
    -- successors 175 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/addr_of_503_complete/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/addr_of_503_complete/final_reg_ack
      -- 
    final_reg_ack_11566_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_503_final_reg_ack_0, ack => cp_elements(189)); -- 
    -- CP-element group 190 join  fork  transition  bypass 
    -- predecessors 194 196 
    -- successors 191 197 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_active_
      -- 
    cpelement_group_190 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(194);
      predecessors(1) <= cp_elements(196);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(190)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(190),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 191 join  fork  transition  place  bypass 
    -- predecessors 190 199 
    -- successors 200 201 
    -- members (13) 
      -- 	branch_block_stmt_323/assign_stmt_511__entry__
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508__exit__
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/assign_stmt_508_trigger_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/assign_stmt_508_active_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/assign_stmt_508_completed_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_completed_
      -- 	branch_block_stmt_323/assign_stmt_511/$entry
      -- 	branch_block_stmt_323/assign_stmt_511/assign_stmt_511_trigger_
      -- 	branch_block_stmt_323/assign_stmt_511/assign_stmt_511_active_
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_510_trigger_
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_510_active_
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_510_completed_
      -- 
    cpelement_group_191 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(190);
      predecessors(1) <= cp_elements(199);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(191)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(191),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 192 transition  input  output  no-bypass 
    -- predecessors 175 
    -- successors 193 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_address_resized
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_addr_resize/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_plus_offset/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_11584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_base_resize_ack_0, ack => cp_elements(192)); -- 
    sum_rename_req_11588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => ptr_deref_507_root_address_inst_req_0); -- 
    -- CP-element group 193 transition  input  output  no-bypass 
    -- predecessors 192 
    -- successors 194 
    -- members (5) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_root_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_plus_offset/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_word_addrgen/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_word_addrgen/root_register_req
      -- 
    sum_rename_ack_11589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_root_address_inst_ack_0, ack => cp_elements(193)); -- 
    root_register_req_11593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => ptr_deref_507_addr_0_req_0); -- 
    -- CP-element group 194 fork  transition  input  no-bypass 
    -- predecessors 193 
    -- successors 190 195 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_trigger_
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_word_address_calculated
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_word_addrgen/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_word_addrgen/root_register_ack
      -- 
    root_register_ack_11594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_addr_0_ack_0, ack => cp_elements(194)); -- 
    -- CP-element group 195 transition  output  bypass 
    -- predecessors 194 
    -- successors 196 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/word_access/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/word_access/word_access_0/rr
      -- 
    cp_elements(195) <= cp_elements(194);
    rr_11604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => ptr_deref_507_load_0_req_0); -- 
    -- CP-element group 196 transition  input  no-bypass 
    -- predecessors 195 
    -- successors 190 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/word_access/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_request/word_access/word_access_0/ra
      -- 
    ra_11605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_load_0_ack_0, ack => cp_elements(196)); -- 
    -- CP-element group 197 transition  output  bypass 
    -- predecessors 190 
    -- successors 198 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/word_access/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/word_access/word_access_0/cr
      -- 
    cp_elements(197) <= cp_elements(190);
    cr_11615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => ptr_deref_507_load_0_req_1); -- 
    -- CP-element group 198 transition  input  output  no-bypass 
    -- predecessors 197 
    -- successors 199 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/word_access/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/merge_req
      -- 
    ca_11616_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_load_0_ack_1, ack => cp_elements(198)); -- 
    merge_req_11617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => ptr_deref_507_gather_scatter_req_0); -- 
    -- CP-element group 199 transition  input  no-bypass 
    -- predecessors 198 
    -- successors 191 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/$exit
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508/ptr_deref_507_complete/merge_ack
      -- 
    merge_ack_11618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_gather_scatter_ack_0, ack => cp_elements(199)); -- 
    -- CP-element group 200 join  fork  transition  place  no-bypass 
    -- predecessors 191 202 
    -- successors 205 207 
    -- members (9) 
      -- 	branch_block_stmt_323/assign_stmt_511__exit__
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523__entry__
      -- 	branch_block_stmt_323/assign_stmt_511/$exit
      -- 	branch_block_stmt_323/assign_stmt_511/assign_stmt_511_completed_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/$entry
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_trigger_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/simple_obj_ref_513_trigger_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/simple_obj_ref_513_active_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/simple_obj_ref_513_completed_
      -- 
    cpelement_group_200 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(191);
      predecessors(1) <= cp_elements(202);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(200)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(200),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 201 fork  transition  bypass 
    -- predecessors 191 
    -- successors 202 203 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_509_trigger_
      -- 
    cp_elements(201) <= cp_elements(191);
    -- CP-element group 202 join  transition  no-bypass 
    -- predecessors 201 204 
    -- successors 200 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_509_active_
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_509_completed_
      -- 
    cpelement_group_202 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(201);
      predecessors(1) <= cp_elements(204);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(202)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(202),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 203 transition  output  bypass 
    -- predecessors 201 
    -- successors 204 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_509_complete/$entry
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_509_complete/pipe_wreq
      -- 
    cp_elements(203) <= cp_elements(201);
    pipe_wreq_11634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => simple_obj_ref_509_inst_req_0); -- 
    -- CP-element group 204 transition  input  no-bypass 
    -- predecessors 203 
    -- successors 202 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_509_complete/$exit
      -- 	branch_block_stmt_323/assign_stmt_511/simple_obj_ref_509_complete/pipe_wack
      -- 
    pipe_wack_11635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_509_inst_ack_0, ack => cp_elements(204)); -- 
    -- CP-element group 205 join  fork  transition  bypass 
    -- predecessors 200 208 
    -- successors 206 209 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_active_
      -- 
    cpelement_group_205 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(200);
      predecessors(1) <= cp_elements(208);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(205)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(205),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 206 join  fork  transition  no-bypass 
    -- predecessors 205 210 
    -- successors 211 213 
    -- members (8) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/assign_stmt_517_trigger_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/assign_stmt_517_active_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/assign_stmt_517_completed_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_completed_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_trigger_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/simple_obj_ref_519_trigger_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/simple_obj_ref_519_active_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/simple_obj_ref_519_completed_
      -- 
    cpelement_group_206 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(205);
      predecessors(1) <= cp_elements(210);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(206)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(206),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 207 transition  output  bypass 
    -- predecessors 200 
    -- successors 208 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Sample/rr
      -- 
    cp_elements(207) <= cp_elements(200);
    rr_11651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => binary_516_inst_req_0); -- 
    -- CP-element group 208 transition  input  no-bypass 
    -- predecessors 207 
    -- successors 205 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Sample/ra
      -- 
    ra_11652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_516_inst_ack_0, ack => cp_elements(208)); -- 
    -- CP-element group 209 transition  output  bypass 
    -- predecessors 205 
    -- successors 210 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Update/cr
      -- 
    cp_elements(209) <= cp_elements(205);
    cr_11656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => binary_516_inst_req_1); -- 
    -- CP-element group 210 transition  input  no-bypass 
    -- predecessors 209 
    -- successors 206 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_516_complete_Update/ca
      -- 
    ca_11657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_516_inst_ack_1, ack => cp_elements(210)); -- 
    -- CP-element group 211 join  fork  transition  bypass 
    -- predecessors 206 214 
    -- successors 212 215 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_active_
      -- 
    cpelement_group_211 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(206);
      predecessors(1) <= cp_elements(214);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(211)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(211),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 212 branch  join  transition  place  no-bypass 
    -- predecessors 211 216 
    -- successors 217 220 
    -- members (7) 
      -- 	branch_block_stmt_323/if_stmt_524__entry__
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523__exit__
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/$exit
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/assign_stmt_523_trigger_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/assign_stmt_523_active_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/assign_stmt_523_completed_
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_completed_
      -- 
    cpelement_group_212 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(211);
      predecessors(1) <= cp_elements(216);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(212)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(212),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 213 transition  output  bypass 
    -- predecessors 206 
    -- successors 214 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Sample/rr
      -- 
    cp_elements(213) <= cp_elements(206);
    rr_11670_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => binary_522_inst_req_0); -- 
    -- CP-element group 214 transition  input  no-bypass 
    -- predecessors 213 
    -- successors 211 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Sample/ra
      -- 
    ra_11671_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_522_inst_ack_0, ack => cp_elements(214)); -- 
    -- CP-element group 215 transition  output  bypass 
    -- predecessors 211 
    -- successors 216 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Update/cr
      -- 
    cp_elements(215) <= cp_elements(211);
    cr_11675_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(215), ack => binary_522_inst_req_1); -- 
    -- CP-element group 216 transition  input  no-bypass 
    -- predecessors 215 
    -- successors 212 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_517_to_assign_stmt_523/binary_522_complete_Update/ca
      -- 
    ca_11676_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_522_inst_ack_1, ack => cp_elements(216)); -- 
    -- CP-element group 217 transition  bypass 
    -- predecessors 212 
    -- successors 218 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_524_dead_link/$entry
      -- 
    cp_elements(217) <= cp_elements(212);
    -- CP-element group 218 transition  dead  bypass 
    -- predecessors 217 
    -- successors 219 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_524_dead_link/dead_transition
      -- 
    cp_elements(218) <= false;
    -- CP-element group 219 transition  place  bypass 
    -- predecessors 218 
    -- successors 283 
    -- members (4) 
      -- 	branch_block_stmt_323/if_stmt_524__exit__
      -- 	branch_block_stmt_323/merge_stmt_530__entry__
      -- 	branch_block_stmt_323/merge_stmt_530_dead_link/$entry
      -- 	branch_block_stmt_323/if_stmt_524_dead_link/$exit
      -- 
    cp_elements(219) <= cp_elements(218);
    -- CP-element group 220 transition  output  bypass 
    -- predecessors 212 
    -- successors 221 
    -- members (3) 
      -- 	branch_block_stmt_323/if_stmt_524_eval_test/$entry
      -- 	branch_block_stmt_323/if_stmt_524_eval_test/$exit
      -- 	branch_block_stmt_323/if_stmt_524_eval_test/branch_req
      -- 
    cp_elements(220) <= cp_elements(212);
    branch_req_11684_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(220), ack => if_stmt_524_branch_req_0); -- 
    -- CP-element group 221 branch  place  bypass 
    -- predecessors 220 
    -- successors 222 224 
    -- members (1) 
      -- 	branch_block_stmt_323/simple_obj_ref_525_place
      -- 
    cp_elements(221) <= cp_elements(220);
    -- CP-element group 222 transition  bypass 
    -- predecessors 221 
    -- successors 223 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_524_if_link/$entry
      -- 
    cp_elements(222) <= cp_elements(221);
    -- CP-element group 223 transition  place  input  no-bypass 
    -- predecessors 222 
    -- successors 7 
    -- members (9) 
      -- 	branch_block_stmt_323/bb_12_xx_x_crit_edgex_xi4_PhiReq/$entry
      -- 	branch_block_stmt_323/merge_stmt_530_PhiAck/$entry
      -- 	branch_block_stmt_323/merge_stmt_530_PhiAck/$exit
      -- 	branch_block_stmt_323/bb_12_xx_x_crit_edgex_xi4_PhiReq/$exit
      -- 	branch_block_stmt_323/merge_stmt_530_PhiReqMerge
      -- 	branch_block_stmt_323/if_stmt_524_if_link/$exit
      -- 	branch_block_stmt_323/if_stmt_524_if_link/if_choice_transition
      -- 	branch_block_stmt_323/bb_12_xx_x_crit_edgex_xi4
      -- 	branch_block_stmt_323/merge_stmt_530_PhiAck/dummy
      -- 
    if_choice_transition_11689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_524_branch_ack_1, ack => cp_elements(223)); -- 
    -- CP-element group 224 transition  bypass 
    -- predecessors 221 
    -- successors 225 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_524_else_link/$entry
      -- 
    cp_elements(224) <= cp_elements(221);
    -- CP-element group 225 transition  place  input  output  no-bypass 
    -- predecessors 224 
    -- successors 279 
    -- members (8) 
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/$entry
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/req
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/$entry
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/$entry
      -- 	branch_block_stmt_323/if_stmt_524_else_link/$exit
      -- 	branch_block_stmt_323/if_stmt_524_else_link/else_choice_transition
      -- 	branch_block_stmt_323/bb_12_bb_12
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/$entry
      -- 
    else_choice_transition_11693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_524_branch_ack_0, ack => cp_elements(225)); -- 
    req_12034_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => type_cast_497_inst_req_0); -- 
    -- CP-element group 226 join  fork  transition  bypass 
    -- predecessors 7 229 
    -- successors 227 230 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_active_
      -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(7);
      predecessors(1) <= cp_elements(229);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(226)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 227 join  fork  transition  bypass 
    -- predecessors 226 231 
    -- successors 232 234 
    -- members (8) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/assign_stmt_536_trigger_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/assign_stmt_536_active_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/assign_stmt_536_completed_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_completed_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_trigger_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/simple_obj_ref_538_trigger_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/simple_obj_ref_538_active_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/simple_obj_ref_538_completed_
      -- 
    cpelement_group_227 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(226);
      predecessors(1) <= cp_elements(231);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(227)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(227),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 228 transition  output  bypass 
    -- predecessors 7 
    -- successors 229 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Sample/rr
      -- 
    cp_elements(228) <= cp_elements(7);
    rr_11711_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => binary_535_inst_req_0); -- 
    -- CP-element group 229 transition  input  no-bypass 
    -- predecessors 228 
    -- successors 226 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Sample/ra
      -- 
    ra_11712_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_535_inst_ack_0, ack => cp_elements(229)); -- 
    -- CP-element group 230 transition  output  bypass 
    -- predecessors 226 
    -- successors 231 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Update/cr
      -- 
    cp_elements(230) <= cp_elements(226);
    cr_11716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => binary_535_inst_req_1); -- 
    -- CP-element group 231 transition  input  no-bypass 
    -- predecessors 230 
    -- successors 227 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_535_complete_Update/ca
      -- 
    ca_11717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_535_inst_ack_1, ack => cp_elements(231)); -- 
    -- CP-element group 232 join  fork  transition  no-bypass 
    -- predecessors 227 235 
    -- successors 233 236 
    -- members (1) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_active_
      -- 
    cpelement_group_232 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(227);
      predecessors(1) <= cp_elements(235);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(232)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(232),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 233 branch  join  transition  place  no-bypass 
    -- predecessors 232 237 
    -- successors 238 241 
    -- members (7) 
      -- 	branch_block_stmt_323/if_stmt_543__entry__
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542__exit__
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/$exit
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/assign_stmt_542_trigger_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/assign_stmt_542_active_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/assign_stmt_542_completed_
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_completed_
      -- 
    cpelement_group_233 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(232);
      predecessors(1) <= cp_elements(237);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(233)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(233),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 234 transition  output  bypass 
    -- predecessors 227 
    -- successors 235 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Sample/$entry
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Sample/rr
      -- 
    cp_elements(234) <= cp_elements(227);
    rr_11730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => binary_541_inst_req_0); -- 
    -- CP-element group 235 transition  input  no-bypass 
    -- predecessors 234 
    -- successors 232 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Sample/$exit
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Sample/ra
      -- 
    ra_11731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_541_inst_ack_0, ack => cp_elements(235)); -- 
    -- CP-element group 236 transition  output  bypass 
    -- predecessors 232 
    -- successors 237 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Update/$entry
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Update/cr
      -- 
    cp_elements(236) <= cp_elements(232);
    cr_11735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => binary_541_inst_req_1); -- 
    -- CP-element group 237 transition  input  no-bypass 
    -- predecessors 236 
    -- successors 233 
    -- members (2) 
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Update/$exit
      -- 	branch_block_stmt_323/assign_stmt_536_to_assign_stmt_542/binary_541_complete_Update/ca
      -- 
    ca_11736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_541_inst_ack_1, ack => cp_elements(237)); -- 
    -- CP-element group 238 transition  bypass 
    -- predecessors 233 
    -- successors 239 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_543_dead_link/$entry
      -- 
    cp_elements(238) <= cp_elements(233);
    -- CP-element group 239 transition  dead  bypass 
    -- predecessors 238 
    -- successors 240 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_543_dead_link/dead_transition
      -- 
    cp_elements(239) <= false;
    -- CP-element group 240 transition  place  bypass 
    -- predecessors 239 
    -- successors 
    -- members (5) 
      -- 	branch_block_stmt_323/if_stmt_543__exit__
      -- 	$exit
      -- 	branch_block_stmt_323/$exit
      -- 	branch_block_stmt_323/branch_block_stmt_323__exit__
      -- 	branch_block_stmt_323/if_stmt_543_dead_link/$exit
      -- 
    cp_elements(240) <= cp_elements(239);
    -- CP-element group 241 transition  output  bypass 
    -- predecessors 233 
    -- successors 242 
    -- members (3) 
      -- 	branch_block_stmt_323/if_stmt_543_eval_test/$entry
      -- 	branch_block_stmt_323/if_stmt_543_eval_test/$exit
      -- 	branch_block_stmt_323/if_stmt_543_eval_test/branch_req
      -- 
    cp_elements(241) <= cp_elements(233);
    branch_req_11744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => if_stmt_543_branch_req_0); -- 
    -- CP-element group 242 branch  place  bypass 
    -- predecessors 241 
    -- successors 243 245 
    -- members (1) 
      -- 	branch_block_stmt_323/simple_obj_ref_544_place
      -- 
    cp_elements(242) <= cp_elements(241);
    -- CP-element group 243 transition  bypass 
    -- predecessors 242 
    -- successors 244 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_543_if_link/$entry
      -- 
    cp_elements(243) <= cp_elements(242);
    -- CP-element group 244 transition  place  input  output  no-bypass 
    -- predecessors 243 
    -- successors 260 
    -- members (22) 
      -- 	branch_block_stmt_323/merge_stmt_325__exit__
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_req
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/ack
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/req
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xloopexit_bbx_xnph11x_xix_xbackedge_PhiReq/$entry
      -- 	branch_block_stmt_323/if_stmt_543_if_link/$exit
      -- 	branch_block_stmt_323/if_stmt_543_if_link/if_choice_transition
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnph11x_xix_xloopexit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnph11x_xix_xloopexit_PhiReq/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnph11x_xix_xloopexit_PhiReq/$exit
      -- 	branch_block_stmt_323/merge_stmt_325_PhiReqMerge
      -- 	branch_block_stmt_323/merge_stmt_325_PhiAck/$entry
      -- 	branch_block_stmt_323/merge_stmt_325_PhiAck/$exit
      -- 	branch_block_stmt_323/merge_stmt_325_PhiAck/dummy
      -- 
    if_choice_transition_11749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_543_branch_ack_1, ack => cp_elements(244)); -- 
    phi_stmt_397_req_11864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => phi_stmt_397_req_1); -- 
    -- CP-element group 245 transition  bypass 
    -- predecessors 242 
    -- successors 246 
    -- members (1) 
      -- 	branch_block_stmt_323/if_stmt_543_else_link/$entry
      -- 
    cp_elements(245) <= cp_elements(242);
    -- CP-element group 246 transition  place  input  output  no-bypass 
    -- predecessors 245 
    -- successors 275 
    -- members (8) 
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/req
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/$entry
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/$entry
      -- 	branch_block_stmt_323/if_stmt_543_else_link/$exit
      -- 	branch_block_stmt_323/if_stmt_543_else_link/else_choice_transition
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1
      -- 
    else_choice_transition_11753_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_543_branch_ack_0, ack => cp_elements(246)); -- 
    req_12014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => type_cast_487_inst_req_0); -- 
    -- CP-element group 247 transition  input  output  no-bypass 
    -- predecessors 3 
    -- successors 248 
    -- members (6) 
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_req
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/ack
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/type_cast_334/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/phi_stmt_328_sources/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/phi_stmt_328/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xix_xbackedge_bbx_xnph11x_xi_PhiReq/$exit
      -- 
    ack_11792_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_334_inst_ack_0, ack => cp_elements(247)); -- 
    phi_stmt_328_req_11793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(247), ack => phi_stmt_328_req_1); -- 
    -- CP-element group 248 merge  place  bypass 
    -- predecessors 0 247 
    -- successors 249 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_327_PhiReqMerge
      -- 
    cp_elements(248) <= OrReduce(cp_elements(0) & cp_elements(247));
    -- CP-element group 249 transition  bypass 
    -- predecessors 248 
    -- successors 250 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_327_PhiAck/$entry
      -- 
    cp_elements(249) <= cp_elements(248);
    -- CP-element group 250 transition  place  input  output  no-bypass 
    -- predecessors 249 
    -- successors 252 
    -- members (15) 
      -- 	branch_block_stmt_323/merge_stmt_327__exit__
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_req
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/ack
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/req
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/phi_stmt_338/$entry
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/$exit
      -- 	branch_block_stmt_323/bbx_xnph11x_xi_bb_3_PhiReq/$entry
      -- 	branch_block_stmt_323/merge_stmt_327_PhiAck/phi_stmt_328_ack
      -- 	branch_block_stmt_323/merge_stmt_327_PhiAck/$exit
      -- 
    phi_stmt_328_ack_11798_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_328_ack_0, ack => cp_elements(250)); -- 
    phi_stmt_338_req_11828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => phi_stmt_338_req_0); -- 
    -- CP-element group 251 transition  input  output  no-bypass 
    -- predecessors 67 
    -- successors 252 
    -- members (6) 
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_req
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/ack
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/$exit
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/phi_stmt_338_sources/$exit
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/phi_stmt_338/$exit
      -- 	branch_block_stmt_323/bb_3_bb_3_PhiReq/$exit
      -- 
    ack_11812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_344_inst_ack_0, ack => cp_elements(251)); -- 
    phi_stmt_338_req_11813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => phi_stmt_338_req_1); -- 
    -- CP-element group 252 merge  place  bypass 
    -- predecessors 250 251 
    -- successors 253 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_337_PhiReqMerge
      -- 
    cp_elements(252) <= OrReduce(cp_elements(250) & cp_elements(251));
    -- CP-element group 253 transition  bypass 
    -- predecessors 252 
    -- successors 254 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_337_PhiAck/$entry
      -- 
    cp_elements(253) <= cp_elements(252);
    -- CP-element group 254 transition  place  input  no-bypass 
    -- predecessors 253 
    -- successors 8 
    -- members (4) 
      -- 	branch_block_stmt_323/merge_stmt_337__exit__
      -- 	branch_block_stmt_323/assign_stmt_351__entry__
      -- 	branch_block_stmt_323/merge_stmt_337_PhiAck/phi_stmt_338_ack
      -- 	branch_block_stmt_323/merge_stmt_337_PhiAck/$exit
      -- 
    phi_stmt_338_ack_11833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_338_ack_0, ack => cp_elements(254)); -- 
    -- CP-element group 255 transition  dead  bypass 
    -- predecessors 61 
    -- successors 256 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_377_dead_link/dead_transition
      -- 
    cp_elements(255) <= false;
    -- CP-element group 256 transition  bypass 
    -- predecessors 255 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_377_dead_link/$exit
      -- 
    cp_elements(256) <= cp_elements(255);
    -- CP-element group 257 transition  dead  bypass 
    -- predecessors 82 
    -- successors 258 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_396_dead_link/dead_transition
      -- 
    cp_elements(257) <= false;
    -- CP-element group 258 transition  bypass 
    -- predecessors 257 
    -- successors 3 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_396_dead_link/$exit
      -- 
    cp_elements(258) <= cp_elements(257);
    -- CP-element group 259 transition  input  output  no-bypass 
    -- predecessors 88 
    -- successors 260 
    -- members (6) 
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_req
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/ack
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/type_cast_400/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/phi_stmt_397_sources/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/phi_stmt_397/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edge12x_xi_bbx_xnph11x_xix_xbackedge_PhiReq/$exit
      -- 
    ack_11878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_400_inst_ack_0, ack => cp_elements(259)); -- 
    phi_stmt_397_req_11879_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => phi_stmt_397_req_0); -- 
    -- CP-element group 260 merge  place  bypass 
    -- predecessors 244 259 
    -- successors 261 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_396_PhiReqMerge
      -- 
    cp_elements(260) <= OrReduce(cp_elements(244) & cp_elements(259));
    -- CP-element group 261 transition  bypass 
    -- predecessors 260 
    -- successors 262 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_396_PhiAck/$entry
      -- 
    cp_elements(261) <= cp_elements(260);
    -- CP-element group 262 transition  input  no-bypass 
    -- predecessors 261 
    -- successors 3 
    -- members (2) 
      -- 	branch_block_stmt_323/merge_stmt_396_PhiAck/phi_stmt_397_ack
      -- 	branch_block_stmt_323/merge_stmt_396_PhiAck/$exit
      -- 
    phi_stmt_397_ack_11884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_397_ack_0, ack => cp_elements(262)); -- 
    -- CP-element group 263 transition  input  output  no-bypass 
    -- predecessors 169 
    -- successors 264 
    -- members (6) 
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_sources/type_cast_412/ack
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi_bbx_xnphx_xi_PhiReq/phi_stmt_409/phi_stmt_409_req
      -- 
    ack_11921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_412_inst_ack_0, ack => cp_elements(263)); -- 
    phi_stmt_409_req_11922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => phi_stmt_409_req_0); -- 
    -- CP-element group 264 merge  place  bypass 
    -- predecessors 86 263 
    -- successors 265 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_408_PhiReqMerge
      -- 
    cp_elements(264) <= OrReduce(cp_elements(86) & cp_elements(263));
    -- CP-element group 265 transition  bypass 
    -- predecessors 264 
    -- successors 266 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_408_PhiAck/$entry
      -- 
    cp_elements(265) <= cp_elements(264);
    -- CP-element group 266 transition  place  input  output  no-bypass 
    -- predecessors 265 
    -- successors 268 
    -- members (15) 
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/req
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/ack
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_req
      -- 	branch_block_stmt_323/merge_stmt_408_PhiAck/$exit
      -- 	branch_block_stmt_323/merge_stmt_408_PhiAck/phi_stmt_409_ack
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/$entry
      -- 	branch_block_stmt_323/merge_stmt_408__exit__
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/phi_stmt_419/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi_bb_8_PhiReq/$entry
      -- 
    phi_stmt_409_ack_11927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_409_ack_0, ack => cp_elements(266)); -- 
    phi_stmt_419_req_11957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => phi_stmt_419_req_0); -- 
    -- CP-element group 267 transition  input  output  no-bypass 
    -- predecessors 148 
    -- successors 268 
    -- members (6) 
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/$exit
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/$exit
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/$exit
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/$exit
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_sources/type_cast_425/ack
      -- 	branch_block_stmt_323/bb_8_bb_8_PhiReq/phi_stmt_419/phi_stmt_419_req
      -- 
    ack_11941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_425_inst_ack_0, ack => cp_elements(267)); -- 
    phi_stmt_419_req_11942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => phi_stmt_419_req_1); -- 
    -- CP-element group 268 merge  place  bypass 
    -- predecessors 266 267 
    -- successors 269 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_418_PhiReqMerge
      -- 
    cp_elements(268) <= OrReduce(cp_elements(266) & cp_elements(267));
    -- CP-element group 269 transition  bypass 
    -- predecessors 268 
    -- successors 270 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_418_PhiAck/$entry
      -- 
    cp_elements(269) <= cp_elements(268);
    -- CP-element group 270 transition  place  input  no-bypass 
    -- predecessors 269 
    -- successors 89 
    -- members (4) 
      -- 	branch_block_stmt_323/merge_stmt_418_PhiAck/$exit
      -- 	branch_block_stmt_323/merge_stmt_418_PhiAck/phi_stmt_419_ack
      -- 	branch_block_stmt_323/merge_stmt_418__exit__
      -- 	branch_block_stmt_323/assign_stmt_432__entry__
      -- 
    phi_stmt_419_ack_11962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_419_ack_0, ack => cp_elements(270)); -- 
    -- CP-element group 271 transition  dead  bypass 
    -- predecessors 142 
    -- successors 272 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_458_dead_link/dead_transition
      -- 
    cp_elements(271) <= false;
    -- CP-element group 272 transition  bypass 
    -- predecessors 271 
    -- successors 5 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_458_dead_link/$exit
      -- 
    cp_elements(272) <= cp_elements(271);
    -- CP-element group 273 transition  dead  bypass 
    -- predecessors 163 
    -- successors 274 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_477_dead_link/dead_transition
      -- 
    cp_elements(273) <= false;
    -- CP-element group 274 transition  bypass 
    -- predecessors 273 
    -- successors 6 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_477_dead_link/$exit
      -- 
    cp_elements(274) <= cp_elements(273);
    -- CP-element group 275 transition  input  output  no-bypass 
    -- predecessors 246 
    -- successors 276 
    -- members (6) 
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_req
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/phi_stmt_481_sources/type_cast_487/ack
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/phi_stmt_481/$exit
      -- 	branch_block_stmt_323/xx_x_crit_edgex_xi4_bbx_xnphx_xi1_PhiReq/$exit
      -- 
    ack_12015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_487_inst_ack_0, ack => cp_elements(275)); -- 
    phi_stmt_481_req_12016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => phi_stmt_481_req_1); -- 
    -- CP-element group 276 merge  place  bypass 
    -- predecessors 171 275 
    -- successors 277 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_480_PhiReqMerge
      -- 
    cp_elements(276) <= OrReduce(cp_elements(171) & cp_elements(275));
    -- CP-element group 277 transition  bypass 
    -- predecessors 276 
    -- successors 278 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_480_PhiAck/$entry
      -- 
    cp_elements(277) <= cp_elements(276);
    -- CP-element group 278 transition  place  input  output  no-bypass 
    -- predecessors 277 
    -- successors 280 
    -- members (15) 
      -- 	branch_block_stmt_323/merge_stmt_480_PhiAck/phi_stmt_481_ack
      -- 	branch_block_stmt_323/merge_stmt_480_PhiAck/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12
      -- 	branch_block_stmt_323/merge_stmt_480__exit__
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_req
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/ack
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/req
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/phi_stmt_491/$entry
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/$exit
      -- 	branch_block_stmt_323/bbx_xnphx_xi1_bb_12_PhiReq/$entry
      -- 
    phi_stmt_481_ack_12021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_481_ack_0, ack => cp_elements(278)); -- 
    phi_stmt_491_req_12051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(278), ack => phi_stmt_491_req_0); -- 
    -- CP-element group 279 transition  input  output  no-bypass 
    -- predecessors 225 
    -- successors 280 
    -- members (6) 
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/$exit
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_req
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/ack
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/type_cast_497/$exit
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/phi_stmt_491_sources/$exit
      -- 	branch_block_stmt_323/bb_12_bb_12_PhiReq/phi_stmt_491/$exit
      -- 
    ack_12035_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_497_inst_ack_0, ack => cp_elements(279)); -- 
    phi_stmt_491_req_12036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => phi_stmt_491_req_1); -- 
    -- CP-element group 280 merge  place  bypass 
    -- predecessors 278 279 
    -- successors 281 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_490_PhiReqMerge
      -- 
    cp_elements(280) <= OrReduce(cp_elements(278) & cp_elements(279));
    -- CP-element group 281 transition  bypass 
    -- predecessors 280 
    -- successors 282 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_490_PhiAck/$entry
      -- 
    cp_elements(281) <= cp_elements(280);
    -- CP-element group 282 transition  place  input  no-bypass 
    -- predecessors 281 
    -- successors 172 
    -- members (4) 
      -- 	branch_block_stmt_323/assign_stmt_504_to_assign_stmt_508__entry__
      -- 	branch_block_stmt_323/merge_stmt_490__exit__
      -- 	branch_block_stmt_323/merge_stmt_490_PhiAck/$exit
      -- 	branch_block_stmt_323/merge_stmt_490_PhiAck/phi_stmt_491_ack
      -- 
    phi_stmt_491_ack_12056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_491_ack_0, ack => cp_elements(282)); -- 
    -- CP-element group 283 transition  dead  bypass 
    -- predecessors 219 
    -- successors 284 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_530_dead_link/dead_transition
      -- 
    cp_elements(283) <= false;
    -- CP-element group 284 transition  bypass 
    -- predecessors 283 
    -- successors 7 
    -- members (1) 
      -- 	branch_block_stmt_323/merge_stmt_530_dead_link/$exit
      -- 
    cp_elements(284) <= cp_elements(283);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_349_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_349_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_349_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_349_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_349_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_349_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_430_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_430_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_430_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_430_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_430_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_430_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_502_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_502_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_502_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_502_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_502_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_502_root_address : std_logic_vector(8 downto 0);
    signal exitcond10_451 : std_logic_vector(0 downto 0);
    signal exitcond11_523 : std_logic_vector(0 downto 0);
    signal exitcond12_542 : std_logic_vector(0 downto 0);
    signal exitcond19x_xi_389 : std_logic_vector(0 downto 0);
    signal exitcond9_370 : std_logic_vector(0 downto 0);
    signal exitcond_470 : std_logic_vector(0 downto 0);
    signal iNsTr_13_435 : std_logic_vector(31 downto 0);
    signal iNsTr_15_445 : std_logic_vector(31 downto 0);
    signal iNsTr_17_464 : std_logic_vector(31 downto 0);
    signal iNsTr_22_508 : std_logic_vector(31 downto 0);
    signal iNsTr_25_517 : std_logic_vector(31 downto 0);
    signal iNsTr_27_536 : std_logic_vector(31 downto 0);
    signal iNsTr_3_354 : std_logic_vector(31 downto 0);
    signal iNsTr_5_364 : std_logic_vector(31 downto 0);
    signal iNsTr_7_383 : std_logic_vector(31 downto 0);
    signal ptr_deref_356_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_356_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_356_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_356_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_356_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_356_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_437_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_437_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_437_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_437_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_437_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_437_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_507_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_507_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_507_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_507_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_507_word_offset_0 : std_logic_vector(8 downto 0);
    signal scevgep18x_xi_351 : std_logic_vector(31 downto 0);
    signal scevgepx_xi2_504 : std_logic_vector(31 downto 0);
    signal scevgepx_xi_432 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_347_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_347_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_348_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_348_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_428_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_428_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_429_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_429_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_500_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_500_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_501_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_501_scaled : std_logic_vector(8 downto 0);
    signal storemerge12x_xi_491 : std_logic_vector(31 downto 0);
    signal storemerge13x_xi_328 : std_logic_vector(31 downto 0);
    signal storemerge13x_xix_xbe_397 : std_logic_vector(31 downto 0);
    signal storemerge16x_xi_409 : std_logic_vector(31 downto 0);
    signal storemerge24x_xi_419 : std_logic_vector(31 downto 0);
    signal storemerge310x_xi_338 : std_logic_vector(31 downto 0);
    signal storemerge3x_xi_481 : std_logic_vector(31 downto 0);
    signal type_cast_332_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_334_wire : std_logic_vector(31 downto 0);
    signal type_cast_342_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_344_wire : std_logic_vector(31 downto 0);
    signal type_cast_362_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_368_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_381_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_387_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_400_wire : std_logic_vector(31 downto 0);
    signal type_cast_403_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_412_wire : std_logic_vector(31 downto 0);
    signal type_cast_415_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_423_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_425_wire : std_logic_vector(31 downto 0);
    signal type_cast_443_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_449_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_462_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_468_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_485_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_487_wire : std_logic_vector(31 downto 0);
    signal type_cast_495_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_497_wire : std_logic_vector(31 downto 0);
    signal type_cast_515_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_521_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_534_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_540_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_349_offset_scale_factor_0 <= "000010000";
    array_obj_ref_349_offset_scale_factor_1 <= "000000001";
    array_obj_ref_349_resized_base_address <= "000000000";
    array_obj_ref_430_offset_scale_factor_0 <= "000010000";
    array_obj_ref_430_offset_scale_factor_1 <= "000000001";
    array_obj_ref_430_resized_base_address <= "000000000";
    array_obj_ref_502_offset_scale_factor_0 <= "000010000";
    array_obj_ref_502_offset_scale_factor_1 <= "000000001";
    array_obj_ref_502_resized_base_address <= "000000000";
    ptr_deref_356_word_offset_0 <= "000000000";
    ptr_deref_437_word_offset_0 <= "000000000";
    ptr_deref_507_word_offset_0 <= "000000000";
    type_cast_332_wire_constant <= "00000000000000000000000000000000";
    type_cast_342_wire_constant <= "00000000000000000000000000000000";
    type_cast_362_wire_constant <= "00000000000000000000000000000001";
    type_cast_368_wire_constant <= "00000000000000000000000000010000";
    type_cast_381_wire_constant <= "00000000000000000000000000000001";
    type_cast_387_wire_constant <= "00000000000000000000000000010000";
    type_cast_403_wire_constant <= "00000000000000000000000000000000";
    type_cast_415_wire_constant <= "00000000000000000000000000000000";
    type_cast_423_wire_constant <= "00000000000000000000000000000000";
    type_cast_443_wire_constant <= "00000000000000000000000000000001";
    type_cast_449_wire_constant <= "00000000000000000000000000010000";
    type_cast_462_wire_constant <= "00000000000000000000000000000001";
    type_cast_468_wire_constant <= "00000000000000000000000000010000";
    type_cast_485_wire_constant <= "00000000000000000000000000000000";
    type_cast_495_wire_constant <= "00000000000000000000000000000000";
    type_cast_515_wire_constant <= "00000000000000000000000000000001";
    type_cast_521_wire_constant <= "00000000000000000000000000010000";
    type_cast_534_wire_constant <= "00000000000000000000000000000001";
    type_cast_540_wire_constant <= "00000000000000000000000000010000";
    phi_stmt_328: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_332_wire_constant & type_cast_334_wire;
      req <= phi_stmt_328_req_0 & phi_stmt_328_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_328_ack_0,
          idata => idata,
          odata => storemerge13x_xi_328,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_328
    phi_stmt_338: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_342_wire_constant & type_cast_344_wire;
      req <= phi_stmt_338_req_0 & phi_stmt_338_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_338_ack_0,
          idata => idata,
          odata => storemerge310x_xi_338,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_338
    phi_stmt_397: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_400_wire & type_cast_403_wire_constant;
      req <= phi_stmt_397_req_0 & phi_stmt_397_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_397_ack_0,
          idata => idata,
          odata => storemerge13x_xix_xbe_397,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_397
    phi_stmt_409: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_412_wire & type_cast_415_wire_constant;
      req <= phi_stmt_409_req_0 & phi_stmt_409_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_409_ack_0,
          idata => idata,
          odata => storemerge16x_xi_409,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_409
    phi_stmt_419: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_423_wire_constant & type_cast_425_wire;
      req <= phi_stmt_419_req_0 & phi_stmt_419_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_419_ack_0,
          idata => idata,
          odata => storemerge24x_xi_419,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_419
    phi_stmt_481: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_485_wire_constant & type_cast_487_wire;
      req <= phi_stmt_481_req_0 & phi_stmt_481_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_481_ack_0,
          idata => idata,
          odata => storemerge3x_xi_481,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_481
    phi_stmt_491: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_495_wire_constant & type_cast_497_wire;
      req <= phi_stmt_491_req_0 & phi_stmt_491_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_491_ack_0,
          idata => idata,
          odata => storemerge12x_xi_491,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_491
    register_block_0 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_350_final_reg_req_0;
      addr_of_350_final_reg_ack_0 <= ack; 
      addr_of_350_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_349_root_address, dout => scevgep18x_xi_351, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_1 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_431_final_reg_req_0;
      addr_of_431_final_reg_ack_0 <= ack; 
      addr_of_431_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_430_root_address, dout => scevgepx_xi_432, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_2 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_503_final_reg_req_0;
      addr_of_503_final_reg_ack_0 <= ack; 
      addr_of_503_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_502_root_address, dout => scevgepx_xi2_504, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_3 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_349_index_0_resize_req_0;
      array_obj_ref_349_index_0_resize_ack_0 <= ack; 
      array_obj_ref_349_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => storemerge13x_xi_328, dout => simple_obj_ref_347_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_4 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_349_index_1_resize_req_0;
      array_obj_ref_349_index_1_resize_ack_0 <= ack; 
      array_obj_ref_349_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => storemerge310x_xi_338, dout => simple_obj_ref_348_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_5 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_349_offset_inst_req_0;
      array_obj_ref_349_offset_inst_ack_0 <= ack; 
      array_obj_ref_349_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_349_index_partial_sum_1, dout => array_obj_ref_349_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_6 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_430_index_0_resize_req_0;
      array_obj_ref_430_index_0_resize_ack_0 <= ack; 
      array_obj_ref_430_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => storemerge16x_xi_409, dout => simple_obj_ref_428_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_7 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_430_index_1_resize_req_0;
      array_obj_ref_430_index_1_resize_ack_0 <= ack; 
      array_obj_ref_430_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => storemerge24x_xi_419, dout => simple_obj_ref_429_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_8 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_430_offset_inst_req_0;
      array_obj_ref_430_offset_inst_ack_0 <= ack; 
      array_obj_ref_430_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_430_index_partial_sum_1, dout => array_obj_ref_430_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_9 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_502_index_0_resize_req_0;
      array_obj_ref_502_index_0_resize_ack_0 <= ack; 
      array_obj_ref_502_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => storemerge3x_xi_481, dout => simple_obj_ref_500_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_10 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_502_index_1_resize_req_0;
      array_obj_ref_502_index_1_resize_ack_0 <= ack; 
      array_obj_ref_502_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => storemerge12x_xi_491, dout => simple_obj_ref_501_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_11 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_502_offset_inst_req_0;
      array_obj_ref_502_offset_inst_ack_0 <= ack; 
      array_obj_ref_502_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_502_index_partial_sum_1, dout => array_obj_ref_502_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_12 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_356_addr_0_req_0;
      ptr_deref_356_addr_0_ack_0 <= ack; 
      ptr_deref_356_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_356_root_address, dout => ptr_deref_356_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_13 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_356_base_resize_req_0;
      ptr_deref_356_base_resize_ack_0 <= ack; 
      ptr_deref_356_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep18x_xi_351, dout => ptr_deref_356_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_14 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_437_addr_0_req_0;
      ptr_deref_437_addr_0_ack_0 <= ack; 
      ptr_deref_437_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_437_root_address, dout => ptr_deref_437_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_15 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_437_base_resize_req_0;
      ptr_deref_437_base_resize_ack_0 <= ack; 
      ptr_deref_437_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgepx_xi_432, dout => ptr_deref_437_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_16 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_507_addr_0_req_0;
      ptr_deref_507_addr_0_ack_0 <= ack; 
      ptr_deref_507_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_507_root_address, dout => ptr_deref_507_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_17 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_507_base_resize_req_0;
      ptr_deref_507_base_resize_ack_0 <= ack; 
      ptr_deref_507_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgepx_xi2_504, dout => ptr_deref_507_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_18 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_334_inst_req_0;
      type_cast_334_inst_ack_0 <= ack; 
      type_cast_334_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => storemerge13x_xix_xbe_397, dout => type_cast_334_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_19 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_344_inst_req_0;
      type_cast_344_inst_ack_0 <= ack; 
      type_cast_344_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_5_364, dout => type_cast_344_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_20 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_400_inst_req_0;
      type_cast_400_inst_ack_0 <= ack; 
      type_cast_400_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_7_383, dout => type_cast_400_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_21 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_412_inst_req_0;
      type_cast_412_inst_ack_0 <= ack; 
      type_cast_412_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_17_464, dout => type_cast_412_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_22 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_425_inst_req_0;
      type_cast_425_inst_ack_0 <= ack; 
      type_cast_425_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_15_445, dout => type_cast_425_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_23 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_487_inst_req_0;
      type_cast_487_inst_ack_0 <= ack; 
      type_cast_487_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_27_536, dout => type_cast_487_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_24 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_497_inst_req_0;
      type_cast_497_inst_ack_0 <= ack; 
      type_cast_497_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_25_517, dout => type_cast_497_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    array_obj_ref_349_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_349_index_1_rename_ack_0 <= array_obj_ref_349_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_348_resized;
      simple_obj_ref_348_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_349_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_349_root_address_inst_ack_0 <= array_obj_ref_349_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_349_final_offset;
      array_obj_ref_349_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_430_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_430_index_1_rename_ack_0 <= array_obj_ref_430_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_429_resized;
      simple_obj_ref_429_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_430_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_430_root_address_inst_ack_0 <= array_obj_ref_430_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_430_final_offset;
      array_obj_ref_430_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_502_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_502_index_1_rename_ack_0 <= array_obj_ref_502_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_501_resized;
      simple_obj_ref_501_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_502_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_502_root_address_inst_ack_0 <= array_obj_ref_502_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_502_final_offset;
      array_obj_ref_502_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_356_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_356_gather_scatter_ack_0 <= ptr_deref_356_gather_scatter_req_0;
      aggregated_sig <= iNsTr_3_354;
      ptr_deref_356_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_356_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_356_root_address_inst_ack_0 <= ptr_deref_356_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_356_resized_base_address;
      ptr_deref_356_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_437_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_437_gather_scatter_ack_0 <= ptr_deref_437_gather_scatter_req_0;
      aggregated_sig <= iNsTr_13_435;
      ptr_deref_437_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_437_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_437_root_address_inst_ack_0 <= ptr_deref_437_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_437_resized_base_address;
      ptr_deref_437_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_507_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_507_gather_scatter_ack_0 <= ptr_deref_507_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_507_data_0;
      iNsTr_22_508 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_507_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_507_root_address_inst_ack_0 <= ptr_deref_507_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_507_resized_base_address;
      ptr_deref_507_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    if_stmt_371_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_370;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_371_branch_req_0,
          ack0 => if_stmt_371_branch_ack_0,
          ack1 => if_stmt_371_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_390_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond19x_xi_389;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_390_branch_req_0,
          ack0 => if_stmt_390_branch_ack_0,
          ack1 => if_stmt_390_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_452_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond10_451;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_452_branch_req_0,
          ack0 => if_stmt_452_branch_ack_0,
          ack1 => if_stmt_452_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_471_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_470;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_471_branch_req_0,
          ack0 => if_stmt_471_branch_ack_0,
          ack1 => if_stmt_471_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_524_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond11_523;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_524_branch_req_0,
          ack0 => if_stmt_524_branch_ack_0,
          ack1 => if_stmt_524_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_543_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond12_542;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_543_branch_req_0,
          ack0 => if_stmt_543_branch_ack_0,
          ack1 => if_stmt_543_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_430_index_0_scale array_obj_ref_502_index_0_scale array_obj_ref_349_index_0_scale 
    ApIntMul_group_0: Block -- 
      signal data_in: std_logic_vector(26 downto 0);
      signal data_out: std_logic_vector(26 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_428_resized & simple_obj_ref_500_resized & simple_obj_ref_347_resized;
      simple_obj_ref_428_scaled <= data_out(26 downto 18);
      simple_obj_ref_500_scaled <= data_out(17 downto 9);
      simple_obj_ref_347_scaled <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      reqL_unguarded(2) <= array_obj_ref_430_index_0_scale_req_0;
      reqL_unguarded(1) <= array_obj_ref_502_index_0_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_349_index_0_scale_req_0;
      array_obj_ref_430_index_0_scale_ack_0 <= ackL_unguarded(2);
      array_obj_ref_502_index_0_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_349_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= array_obj_ref_430_index_0_scale_req_1;
      reqR_unguarded(1) <= array_obj_ref_502_index_0_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_349_index_0_scale_req_1;
      array_obj_ref_430_index_0_scale_ack_1 <= ackR_unguarded(2);
      array_obj_ref_502_index_0_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_349_index_0_scale_ack_1 <= ackR_unguarded(0);
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000010000",
          constant_width => 9,
          use_constant  => true,
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 3--
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_349_index_sum_1 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_348_scaled & simple_obj_ref_347_scaled;
      array_obj_ref_349_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_349_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_349_index_sum_1_req_1;
      array_obj_ref_349_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_349_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_430_index_sum_1 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_429_scaled & simple_obj_ref_428_scaled;
      array_obj_ref_430_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_430_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_430_index_sum_1_req_1;
      array_obj_ref_430_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_430_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_502_index_sum_1 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_501_scaled & simple_obj_ref_500_scaled;
      array_obj_ref_502_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_502_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_502_index_sum_1_req_1;
      array_obj_ref_502_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_502_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_363_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= storemerge310x_xi_338;
      iNsTr_5_364 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_363_inst_req_0;
      reqR(0) <= binary_363_inst_req_1;
      binary_363_inst_ack_0 <= ackL(0); 
      binary_363_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_369_inst 
    ApIntEq_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_5_364;
      exitcond9_370 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_369_inst_req_0;
      reqR(0) <= binary_369_inst_req_1;
      binary_369_inst_ack_0 <= ackL(0); 
      binary_369_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_382_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= storemerge13x_xi_328;
      iNsTr_7_383 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_382_inst_req_0;
      reqR(0) <= binary_382_inst_req_1;
      binary_382_inst_ack_0 <= ackL(0); 
      binary_382_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_388_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_7_383;
      exitcond19x_xi_389 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_388_inst_req_0;
      reqR(0) <= binary_388_inst_req_1;
      binary_388_inst_ack_0 <= ackL(0); 
      binary_388_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_444_inst 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= storemerge24x_xi_419;
      iNsTr_15_445 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_444_inst_req_0;
      reqR(0) <= binary_444_inst_req_1;
      binary_444_inst_ack_0 <= ackL(0); 
      binary_444_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_450_inst 
    ApIntEq_group_9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_15_445;
      exitcond10_451 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_450_inst_req_0;
      reqR(0) <= binary_450_inst_req_1;
      binary_450_inst_ack_0 <= ackL(0); 
      binary_450_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_463_inst 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= storemerge16x_xi_409;
      iNsTr_17_464 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_463_inst_req_0;
      reqR(0) <= binary_463_inst_req_1;
      binary_463_inst_ack_0 <= ackL(0); 
      binary_463_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_469_inst 
    ApIntEq_group_11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_17_464;
      exitcond_470 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_469_inst_req_0;
      reqR(0) <= binary_469_inst_req_1;
      binary_469_inst_ack_0 <= ackL(0); 
      binary_469_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : binary_516_inst 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= storemerge12x_xi_491;
      iNsTr_25_517 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_516_inst_req_0;
      reqR(0) <= binary_516_inst_req_1;
      binary_516_inst_ack_0 <= ackL(0); 
      binary_516_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_522_inst 
    ApIntEq_group_13: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_25_517;
      exitcond11_523 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_522_inst_req_0;
      reqR(0) <= binary_522_inst_req_1;
      binary_522_inst_ack_0 <= ackL(0); 
      binary_522_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_535_inst 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= storemerge3x_xi_481;
      iNsTr_27_536 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_535_inst_req_0;
      reqR(0) <= binary_535_inst_req_1;
      binary_535_inst_ack_0 <= ackL(0); 
      binary_535_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_541_inst 
    ApIntEq_group_15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_27_536;
      exitcond12_542 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_541_inst_req_0;
      reqR(0) <= binary_541_inst_req_1;
      binary_541_inst_ack_0 <= ackL(0); 
      binary_541_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared load operator group (0) : ptr_deref_507_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_507_load_0_req_0;
      ptr_deref_507_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_507_load_0_req_1;
      ptr_deref_507_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_507_word_address_0;
      ptr_deref_507_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 9,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(8 downto 0),
          mtag => memory_space_2_lr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_356_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(8 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_356_store_0_req_0;
      ptr_deref_356_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_356_store_0_req_1;
      ptr_deref_356_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_356_word_address_0;
      data_in <= ptr_deref_356_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 9,
        data_width => 32,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(8 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_437_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(8 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_437_store_0_req_0;
      ptr_deref_437_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_437_store_0_req_1;
      ptr_deref_437_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_437_word_address_0;
      data_in <= ptr_deref_437_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 9,
        data_width => 32,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(8 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : simple_obj_ref_353_inst simple_obj_ref_434_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      signal req_unguarded, ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      -- 
    begin -- 
      req_unguarded(1) <= simple_obj_ref_353_inst_req_0;
      req_unguarded(0) <= simple_obj_ref_434_inst_req_0;
      simple_obj_ref_353_inst_ack_0 <= ack_unguarded(1);
      simple_obj_ref_434_inst_ack_0 <= ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => req_unguarded,
        ackL => ack_unguarded,
        reqR => req,
        ackR => ack,
        guards => guard_vector); -- 
      iNsTr_3_354 <= data_out(63 downto 32);
      iNsTr_13_435 <= data_out(31 downto 0);
      in_data_pipe_read_0: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 2,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_pipe_read_req(0),
          oack => in_data_pipe_pipe_read_ack(0),
          odata => in_data_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : simple_obj_ref_509_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      signal req_unguarded, ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      req_unguarded(0) <= simple_obj_ref_509_inst_req_0;
      simple_obj_ref_509_inst_ack_0 <= ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => req_unguarded,
        ackL => ack_unguarded,
        reqR => req,
        ackR => ack,
        guards => guard_vector); -- 
      data_in <= iNsTr_22_508;
      result_pipe_write_0: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => result_pipe_pipe_write_req(0),
          oack => result_pipe_pipe_write_ack(0),
          odata => result_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_478_call 
    mmultiply_base_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_478_call_req_0;
      call_stmt_478_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_478_call_req_1;
      call_stmt_478_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => mmultiply_base_call_reqs(0),
          ackR => mmultiply_base_call_acks(0),
          tagR => mmultiply_base_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1, no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => mmultiply_base_return_acks(0), -- cross-over
          ackL => mmultiply_base_return_reqs(0), -- cross-over
          tagL => mmultiply_base_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity mmultiply_base is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(8 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity mmultiply_base;
architecture Default of mmultiply_base is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal mmultiply_base_CP_1311_start: Boolean;
  -- links between control-path and data-path
  signal addr_of_703_final_reg_ack_0 : boolean;
  signal binary_601_inst_req_1 : boolean;
  signal array_obj_ref_696_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_696_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_606_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_606_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_606_index_0_scale_req_0 : boolean;
  signal binary_601_inst_ack_0 : boolean;
  signal array_obj_ref_618_index_0_resize_req_0 : boolean;
  signal array_obj_ref_606_index_sum_1_req_1 : boolean;
  signal array_obj_ref_696_offset_inst_ack_0 : boolean;
  signal array_obj_ref_606_index_0_scale_req_1 : boolean;
  signal array_obj_ref_606_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_708_index_0_scale_req_0 : boolean;
  signal array_obj_ref_630_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_606_offset_inst_req_0 : boolean;
  signal binary_625_inst_ack_1 : boolean;
  signal array_obj_ref_630_index_1_rename_req_0 : boolean;
  signal binary_625_inst_req_0 : boolean;
  signal array_obj_ref_618_root_address_inst_req_0 : boolean;
  signal array_obj_ref_606_offset_inst_ack_0 : boolean;
  signal array_obj_ref_606_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_950_index_1_resize_req_0 : boolean;
  signal array_obj_ref_702_index_sum_1_req_1 : boolean;
  signal binary_613_inst_ack_1 : boolean;
  signal array_obj_ref_708_index_1_resize_req_0 : boolean;
  signal array_obj_ref_696_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_708_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_606_root_address_inst_req_0 : boolean;
  signal array_obj_ref_618_offset_inst_req_0 : boolean;
  signal array_obj_ref_618_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_630_offset_inst_ack_0 : boolean;
  signal array_obj_ref_708_index_1_rename_req_0 : boolean;
  signal array_obj_ref_630_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_630_root_address_inst_req_0 : boolean;
  signal array_obj_ref_606_root_address_inst_ack_0 : boolean;
  signal binary_613_inst_req_0 : boolean;
  signal array_obj_ref_618_index_sum_1_req_1 : boolean;
  signal binary_613_inst_ack_0 : boolean;
  signal array_obj_ref_606_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1046_index_1_rename_req_0 : boolean;
  signal array_obj_ref_702_index_0_resize_req_0 : boolean;
  signal array_obj_ref_630_index_sum_1_req_1 : boolean;
  signal addr_of_607_final_reg_req_0 : boolean;
  signal array_obj_ref_950_root_address_inst_req_0 : boolean;
  signal addr_of_607_final_reg_ack_0 : boolean;
  signal array_obj_ref_696_index_0_scale_req_0 : boolean;
  signal array_obj_ref_630_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_702_index_0_scale_ack_0 : boolean;
  signal addr_of_933_final_reg_ack_0 : boolean;
  signal binary_601_inst_ack_1 : boolean;
  signal addr_of_691_final_reg_ack_0 : boolean;
  signal array_obj_ref_618_index_1_resize_req_0 : boolean;
  signal array_obj_ref_702_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_956_index_0_resize_req_0 : boolean;
  signal array_obj_ref_690_root_address_inst_ack_0 : boolean;
  signal binary_625_inst_req_1 : boolean;
  signal array_obj_ref_606_index_0_resize_req_0 : boolean;
  signal array_obj_ref_618_index_sum_1_req_0 : boolean;
  signal array_obj_ref_702_index_0_scale_req_0 : boolean;
  signal binary_585_inst_ack_0 : boolean;
  signal addr_of_631_final_reg_ack_0 : boolean;
  signal array_obj_ref_696_root_address_inst_req_0 : boolean;
  signal binary_579_inst_req_1 : boolean;
  signal array_obj_ref_630_index_sum_1_ack_1 : boolean;
  signal binary_579_inst_ack_1 : boolean;
  signal array_obj_ref_702_offset_inst_ack_0 : boolean;
  signal binary_585_inst_req_0 : boolean;
  signal array_obj_ref_944_index_0_scale_req_0 : boolean;
  signal array_obj_ref_696_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_618_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_950_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_702_index_0_scale_req_1 : boolean;
  signal array_obj_ref_708_index_0_resize_ack_0 : boolean;
  signal binary_579_inst_ack_0 : boolean;
  signal array_obj_ref_630_index_1_resize_req_0 : boolean;
  signal array_obj_ref_630_offset_inst_req_0 : boolean;
  signal array_obj_ref_618_index_1_rename_req_0 : boolean;
  signal addr_of_951_final_reg_ack_0 : boolean;
  signal array_obj_ref_956_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_630_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_630_root_address_inst_ack_0 : boolean;
  signal binary_601_inst_req_0 : boolean;
  signal array_obj_ref_618_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_630_index_0_resize_req_0 : boolean;
  signal array_obj_ref_702_root_address_inst_req_0 : boolean;
  signal array_obj_ref_708_index_0_scale_ack_1 : boolean;
  signal addr_of_619_final_reg_ack_0 : boolean;
  signal binary_625_inst_ack_0 : boolean;
  signal array_obj_ref_630_index_sum_1_req_0 : boolean;
  signal array_obj_ref_956_index_0_scale_req_0 : boolean;
  signal addr_of_631_final_reg_req_0 : boolean;
  signal array_obj_ref_696_index_0_resize_ack_0 : boolean;
  signal addr_of_619_final_reg_req_0 : boolean;
  signal array_obj_ref_606_index_0_resize_ack_0 : boolean;
  signal addr_of_933_final_reg_req_0 : boolean;
  signal binary_585_inst_req_1 : boolean;
  signal binary_613_inst_req_1 : boolean;
  signal binary_585_inst_ack_1 : boolean;
  signal array_obj_ref_630_index_sum_1_ack_0 : boolean;
  signal binary_579_inst_req_0 : boolean;
  signal array_obj_ref_696_index_0_scale_req_1 : boolean;
  signal addr_of_691_final_reg_req_0 : boolean;
  signal array_obj_ref_618_offset_inst_ack_0 : boolean;
  signal array_obj_ref_606_index_1_rename_req_0 : boolean;
  signal array_obj_ref_606_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_690_root_address_inst_req_0 : boolean;
  signal array_obj_ref_606_index_sum_1_req_0 : boolean;
  signal array_obj_ref_606_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_630_index_0_scale_req_1 : boolean;
  signal array_obj_ref_956_index_0_scale_ack_1 : boolean;
  signal binary_573_inst_ack_1 : boolean;
  signal binary_573_inst_req_1 : boolean;
  signal array_obj_ref_618_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_702_index_1_resize_ack_0 : boolean;
  signal binary_573_inst_ack_0 : boolean;
  signal binary_573_inst_req_0 : boolean;
  signal array_obj_ref_702_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_618_index_0_scale_req_1 : boolean;
  signal array_obj_ref_708_index_0_resize_req_0 : boolean;
  signal array_obj_ref_618_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_618_index_0_scale_req_0 : boolean;
  signal binary_567_inst_ack_1 : boolean;
  signal binary_567_inst_req_1 : boolean;
  signal array_obj_ref_630_index_0_scale_ack_0 : boolean;
  signal binary_567_inst_ack_0 : boolean;
  signal array_obj_ref_618_index_1_rename_ack_0 : boolean;
  signal binary_567_inst_req_0 : boolean;
  signal array_obj_ref_702_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_696_offset_inst_req_0 : boolean;
  signal array_obj_ref_950_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_618_root_address_inst_ack_0 : boolean;
  signal phi_stmt_764_req_0 : boolean;
  signal array_obj_ref_690_offset_inst_ack_0 : boolean;
  signal array_obj_ref_630_index_0_scale_req_0 : boolean;
  signal array_obj_ref_618_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_702_offset_inst_req_0 : boolean;
  signal addr_of_697_final_reg_req_0 : boolean;
  signal array_obj_ref_690_index_0_resize_req_0 : boolean;
  signal array_obj_ref_690_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_690_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_932_offset_inst_ack_0 : boolean;
  signal array_obj_ref_708_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_708_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1052_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_932_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_690_index_1_resize_req_0 : boolean;
  signal array_obj_ref_714_index_sum_1_req_1 : boolean;
  signal array_obj_ref_714_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_690_index_0_scale_req_0 : boolean;
  signal array_obj_ref_956_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_690_index_0_scale_ack_0 : boolean;
  signal addr_of_945_final_reg_req_0 : boolean;
  signal array_obj_ref_708_index_1_rename_ack_0 : boolean;
  signal binary_721_inst_req_0 : boolean;
  signal array_obj_ref_950_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_702_index_1_resize_req_0 : boolean;
  signal array_obj_ref_714_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_696_index_1_resize_req_0 : boolean;
  signal array_obj_ref_690_index_0_scale_req_1 : boolean;
  signal array_obj_ref_944_index_0_resize_req_0 : boolean;
  signal array_obj_ref_702_index_sum_1_req_0 : boolean;
  signal array_obj_ref_932_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_714_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1052_index_0_scale_req_0 : boolean;
  signal addr_of_957_final_reg_req_0 : boolean;
  signal binary_721_inst_ack_0 : boolean;
  signal array_obj_ref_702_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_944_index_0_scale_ack_0 : boolean;
  signal binary_727_inst_req_0 : boolean;
  signal array_obj_ref_932_index_0_scale_ack_1 : boolean;
  signal binary_727_inst_ack_0 : boolean;
  signal array_obj_ref_932_offset_inst_req_0 : boolean;
  signal array_obj_ref_708_offset_inst_ack_0 : boolean;
  signal array_obj_ref_950_index_0_resize_req_0 : boolean;
  signal array_obj_ref_696_index_1_resize_ack_0 : boolean;
  signal binary_721_inst_req_1 : boolean;
  signal array_obj_ref_702_root_address_inst_ack_0 : boolean;
  signal binary_721_inst_ack_1 : boolean;
  signal array_obj_ref_1046_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_708_index_sum_1_req_0 : boolean;
  signal addr_of_697_final_reg_ack_0 : boolean;
  signal array_obj_ref_708_index_0_scale_req_1 : boolean;
  signal addr_of_703_final_reg_req_0 : boolean;
  signal array_obj_ref_690_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_950_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_702_index_sum_1_ack_0 : boolean;
  signal binary_1143_inst_ack_1 : boolean;
  signal array_obj_ref_932_index_0_scale_req_1 : boolean;
  signal binary_727_inst_req_1 : boolean;
  signal array_obj_ref_1046_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_962_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_932_index_0_scale_ack_0 : boolean;
  signal binary_727_inst_ack_1 : boolean;
  signal array_obj_ref_932_index_0_scale_req_0 : boolean;
  signal array_obj_ref_684_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_956_root_address_inst_req_0 : boolean;
  signal array_obj_ref_932_root_address_inst_req_0 : boolean;
  signal array_obj_ref_636_index_0_resize_req_0 : boolean;
  signal array_obj_ref_636_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_636_index_0_scale_req_0 : boolean;
  signal array_obj_ref_636_index_0_scale_ack_0 : boolean;
  signal addr_of_685_final_reg_ack_0 : boolean;
  signal array_obj_ref_636_index_0_scale_req_1 : boolean;
  signal addr_of_685_final_reg_req_0 : boolean;
  signal array_obj_ref_636_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_932_index_1_resize_req_0 : boolean;
  signal array_obj_ref_684_root_address_inst_req_0 : boolean;
  signal array_obj_ref_956_index_sum_1_req_1 : boolean;
  signal array_obj_ref_636_index_1_resize_req_0 : boolean;
  signal array_obj_ref_636_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_684_offset_inst_ack_0 : boolean;
  signal array_obj_ref_636_index_1_rename_req_0 : boolean;
  signal array_obj_ref_684_offset_inst_req_0 : boolean;
  signal array_obj_ref_636_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_956_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_684_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_636_index_sum_1_req_0 : boolean;
  signal array_obj_ref_684_index_sum_1_req_1 : boolean;
  signal array_obj_ref_636_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_684_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_636_index_sum_1_req_1 : boolean;
  signal array_obj_ref_684_index_sum_1_req_0 : boolean;
  signal array_obj_ref_636_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_636_offset_inst_req_0 : boolean;
  signal array_obj_ref_636_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1046_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1052_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_684_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_636_root_address_inst_req_0 : boolean;
  signal array_obj_ref_684_index_1_rename_req_0 : boolean;
  signal array_obj_ref_636_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_714_index_1_rename_ack_0 : boolean;
  signal addr_of_637_final_reg_req_0 : boolean;
  signal addr_of_637_final_reg_ack_0 : boolean;
  signal array_obj_ref_714_root_address_inst_req_0 : boolean;
  signal array_obj_ref_684_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_684_index_1_resize_req_0 : boolean;
  signal array_obj_ref_696_index_sum_1_req_1 : boolean;
  signal array_obj_ref_696_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_708_offset_inst_req_0 : boolean;
  signal array_obj_ref_1052_index_sum_1_req_0 : boolean;
  signal array_obj_ref_684_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_684_index_0_scale_req_1 : boolean;
  signal addr_of_945_final_reg_ack_0 : boolean;
  signal array_obj_ref_932_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_684_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_642_index_0_resize_req_0 : boolean;
  signal array_obj_ref_684_index_0_scale_req_0 : boolean;
  signal array_obj_ref_642_index_0_resize_ack_0 : boolean;
  signal addr_of_957_final_reg_ack_0 : boolean;
  signal array_obj_ref_642_index_0_scale_req_0 : boolean;
  signal array_obj_ref_642_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_684_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_642_index_0_scale_req_1 : boolean;
  signal array_obj_ref_684_index_0_resize_req_0 : boolean;
  signal array_obj_ref_642_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_714_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_714_index_0_resize_req_0 : boolean;
  signal array_obj_ref_642_index_1_resize_req_0 : boolean;
  signal array_obj_ref_642_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_714_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1052_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_642_index_1_rename_req_0 : boolean;
  signal array_obj_ref_642_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_932_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_642_index_sum_1_req_0 : boolean;
  signal array_obj_ref_642_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_642_index_sum_1_req_1 : boolean;
  signal array_obj_ref_642_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_642_offset_inst_req_0 : boolean;
  signal array_obj_ref_642_offset_inst_ack_0 : boolean;
  signal array_obj_ref_642_root_address_inst_req_0 : boolean;
  signal array_obj_ref_642_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_714_index_1_rename_req_0 : boolean;
  signal addr_of_679_final_reg_ack_0 : boolean;
  signal addr_of_643_final_reg_req_0 : boolean;
  signal addr_of_679_final_reg_req_0 : boolean;
  signal addr_of_643_final_reg_ack_0 : boolean;
  signal array_obj_ref_708_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_708_root_address_inst_req_0 : boolean;
  signal array_obj_ref_932_index_sum_1_req_1 : boolean;
  signal array_obj_ref_696_index_sum_1_req_0 : boolean;
  signal array_obj_ref_678_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_678_root_address_inst_req_0 : boolean;
  signal array_obj_ref_708_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_678_offset_inst_ack_0 : boolean;
  signal array_obj_ref_678_offset_inst_req_0 : boolean;
  signal array_obj_ref_678_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_678_index_sum_1_req_1 : boolean;
  signal array_obj_ref_678_index_sum_1_ack_0 : boolean;
  signal addr_of_951_final_reg_req_0 : boolean;
  signal array_obj_ref_678_index_sum_1_req_0 : boolean;
  signal array_obj_ref_648_index_0_resize_req_0 : boolean;
  signal array_obj_ref_648_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_714_index_1_resize_req_0 : boolean;
  signal array_obj_ref_648_index_0_scale_req_0 : boolean;
  signal array_obj_ref_678_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_648_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_678_index_1_rename_req_0 : boolean;
  signal array_obj_ref_648_index_0_scale_req_1 : boolean;
  signal array_obj_ref_648_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_678_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_678_index_1_resize_req_0 : boolean;
  signal array_obj_ref_956_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_648_index_1_resize_req_0 : boolean;
  signal array_obj_ref_648_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_648_index_1_rename_req_0 : boolean;
  signal array_obj_ref_648_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_714_offset_inst_ack_0 : boolean;
  signal array_obj_ref_956_offset_inst_ack_0 : boolean;
  signal array_obj_ref_648_index_sum_1_req_0 : boolean;
  signal array_obj_ref_648_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_678_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_648_index_sum_1_req_1 : boolean;
  signal array_obj_ref_678_index_0_scale_req_1 : boolean;
  signal array_obj_ref_648_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_678_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_648_offset_inst_req_0 : boolean;
  signal array_obj_ref_678_index_0_scale_req_0 : boolean;
  signal array_obj_ref_648_offset_inst_ack_0 : boolean;
  signal array_obj_ref_932_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_714_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_648_root_address_inst_req_0 : boolean;
  signal array_obj_ref_648_root_address_inst_ack_0 : boolean;
  signal addr_of_715_final_reg_ack_0 : boolean;
  signal array_obj_ref_678_index_0_resize_ack_0 : boolean;
  signal addr_of_649_final_reg_req_0 : boolean;
  signal array_obj_ref_678_index_0_resize_req_0 : boolean;
  signal addr_of_649_final_reg_ack_0 : boolean;
  signal array_obj_ref_696_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_708_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1052_index_sum_1_req_1 : boolean;
  signal array_obj_ref_956_offset_inst_req_0 : boolean;
  signal array_obj_ref_956_index_0_scale_ack_0 : boolean;
  signal binary_655_inst_req_0 : boolean;
  signal binary_655_inst_ack_0 : boolean;
  signal binary_655_inst_req_1 : boolean;
  signal binary_655_inst_ack_1 : boolean;
  signal array_obj_ref_714_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_944_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_696_index_1_rename_req_0 : boolean;
  signal addr_of_709_final_reg_ack_0 : boolean;
  signal array_obj_ref_1052_index_1_resize_ack_0 : boolean;
  signal addr_of_673_final_reg_ack_0 : boolean;
  signal addr_of_673_final_reg_req_0 : boolean;
  signal array_obj_ref_672_root_address_inst_ack_0 : boolean;
  signal addr_of_709_final_reg_req_0 : boolean;
  signal array_obj_ref_714_index_0_scale_req_1 : boolean;
  signal array_obj_ref_672_root_address_inst_req_0 : boolean;
  signal array_obj_ref_660_index_0_resize_req_0 : boolean;
  signal array_obj_ref_660_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_932_index_1_rename_req_0 : boolean;
  signal addr_of_715_final_reg_req_0 : boolean;
  signal array_obj_ref_660_index_0_scale_req_0 : boolean;
  signal array_obj_ref_672_offset_inst_ack_0 : boolean;
  signal array_obj_ref_660_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_672_offset_inst_req_0 : boolean;
  signal array_obj_ref_660_index_0_scale_req_1 : boolean;
  signal array_obj_ref_672_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_660_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_714_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_672_index_sum_1_req_1 : boolean;
  signal array_obj_ref_672_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_672_index_sum_1_req_0 : boolean;
  signal array_obj_ref_660_index_1_resize_req_0 : boolean;
  signal array_obj_ref_672_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_660_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_672_index_1_rename_req_0 : boolean;
  signal array_obj_ref_660_index_1_rename_req_0 : boolean;
  signal array_obj_ref_660_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_714_offset_inst_req_0 : boolean;
  signal array_obj_ref_950_index_0_scale_req_1 : boolean;
  signal array_obj_ref_932_index_sum_1_req_0 : boolean;
  signal array_obj_ref_714_index_0_scale_req_0 : boolean;
  signal array_obj_ref_660_index_sum_1_req_0 : boolean;
  signal array_obj_ref_672_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_660_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_672_index_1_resize_req_0 : boolean;
  signal array_obj_ref_660_index_sum_1_req_1 : boolean;
  signal array_obj_ref_660_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_660_offset_inst_req_0 : boolean;
  signal array_obj_ref_660_offset_inst_ack_0 : boolean;
  signal array_obj_ref_660_root_address_inst_req_0 : boolean;
  signal array_obj_ref_660_root_address_inst_ack_0 : boolean;
  signal addr_of_661_final_reg_req_0 : boolean;
  signal addr_of_661_final_reg_ack_0 : boolean;
  signal array_obj_ref_690_offset_inst_req_0 : boolean;
  signal array_obj_ref_696_index_0_resize_req_0 : boolean;
  signal array_obj_ref_690_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_690_index_sum_1_req_1 : boolean;
  signal array_obj_ref_690_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_672_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_672_index_0_scale_req_1 : boolean;
  signal array_obj_ref_690_index_sum_1_req_0 : boolean;
  signal array_obj_ref_672_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_672_index_0_scale_req_0 : boolean;
  signal array_obj_ref_672_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_672_index_0_resize_req_0 : boolean;
  signal array_obj_ref_690_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_690_index_1_rename_req_0 : boolean;
  signal array_obj_ref_666_index_0_resize_req_0 : boolean;
  signal array_obj_ref_666_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_666_index_0_scale_req_0 : boolean;
  signal array_obj_ref_666_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_666_index_0_scale_req_1 : boolean;
  signal array_obj_ref_666_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_702_index_1_rename_req_0 : boolean;
  signal array_obj_ref_944_index_0_scale_req_1 : boolean;
  signal array_obj_ref_944_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1046_index_sum_1_req_1 : boolean;
  signal array_obj_ref_666_index_1_resize_req_0 : boolean;
  signal array_obj_ref_666_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_666_index_1_rename_req_0 : boolean;
  signal array_obj_ref_666_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_666_index_sum_1_req_0 : boolean;
  signal array_obj_ref_666_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_666_index_sum_1_req_1 : boolean;
  signal array_obj_ref_666_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_666_offset_inst_req_0 : boolean;
  signal array_obj_ref_666_offset_inst_ack_0 : boolean;
  signal array_obj_ref_950_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_666_root_address_inst_req_0 : boolean;
  signal array_obj_ref_666_root_address_inst_ack_0 : boolean;
  signal addr_of_667_final_reg_req_0 : boolean;
  signal addr_of_667_final_reg_ack_0 : boolean;
  signal array_obj_ref_932_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1046_index_1_resize_req_0 : boolean;
  signal array_obj_ref_932_index_0_resize_req_0 : boolean;
  signal array_obj_ref_962_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_962_index_0_scale_req_1 : boolean;
  signal array_obj_ref_956_index_1_rename_ack_0 : boolean;
  signal binary_733_inst_req_0 : boolean;
  signal binary_733_inst_ack_0 : boolean;
  signal binary_733_inst_req_1 : boolean;
  signal binary_733_inst_ack_1 : boolean;
  signal array_obj_ref_962_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_962_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_962_index_0_scale_req_0 : boolean;
  signal array_obj_ref_962_index_0_resize_req_0 : boolean;
  signal array_obj_ref_950_index_0_scale_req_0 : boolean;
  signal array_obj_ref_956_index_1_rename_req_0 : boolean;
  signal binary_739_inst_req_0 : boolean;
  signal binary_739_inst_ack_0 : boolean;
  signal binary_739_inst_req_1 : boolean;
  signal binary_739_inst_ack_1 : boolean;
  signal addr_of_927_final_reg_ack_0 : boolean;
  signal addr_of_927_final_reg_req_0 : boolean;
  signal array_obj_ref_926_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_944_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1052_index_0_resize_req_0 : boolean;
  signal array_obj_ref_926_root_address_inst_req_0 : boolean;
  signal binary_867_inst_req_0 : boolean;
  signal binary_867_inst_ack_0 : boolean;
  signal binary_867_inst_req_1 : boolean;
  signal array_obj_ref_926_offset_inst_ack_0 : boolean;
  signal binary_867_inst_ack_1 : boolean;
  signal array_obj_ref_956_index_sum_1_req_0 : boolean;
  signal array_obj_ref_962_index_1_resize_req_0 : boolean;
  signal array_obj_ref_926_offset_inst_req_0 : boolean;
  signal array_obj_ref_926_index_sum_1_ack_1 : boolean;
  signal addr_of_939_final_reg_ack_0 : boolean;
  signal array_obj_ref_926_index_sum_1_req_1 : boolean;
  signal array_obj_ref_926_index_sum_1_ack_0 : boolean;
  signal ptr_deref_1125_addr_0_req_0 : boolean;
  signal array_obj_ref_1046_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_926_index_sum_1_req_0 : boolean;
  signal array_obj_ref_926_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_926_index_1_rename_req_0 : boolean;
  signal array_obj_ref_950_offset_inst_ack_0 : boolean;
  signal addr_of_939_final_reg_req_0 : boolean;
  signal array_obj_ref_944_root_address_inst_req_0 : boolean;
  signal array_obj_ref_926_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_872_index_0_resize_req_0 : boolean;
  signal array_obj_ref_926_index_1_resize_req_0 : boolean;
  signal array_obj_ref_872_index_0_resize_ack_0 : boolean;
  signal binary_1148_inst_req_0 : boolean;
  signal array_obj_ref_872_index_0_scale_req_0 : boolean;
  signal array_obj_ref_872_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_872_index_0_scale_req_1 : boolean;
  signal array_obj_ref_872_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_938_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_938_root_address_inst_req_0 : boolean;
  signal array_obj_ref_926_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_950_offset_inst_req_0 : boolean;
  signal array_obj_ref_938_offset_inst_ack_0 : boolean;
  signal array_obj_ref_956_index_0_scale_req_1 : boolean;
  signal array_obj_ref_938_offset_inst_req_0 : boolean;
  signal array_obj_ref_926_index_0_scale_req_1 : boolean;
  signal array_obj_ref_872_index_1_resize_req_0 : boolean;
  signal array_obj_ref_926_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_872_index_1_resize_ack_0 : boolean;
  signal ptr_deref_1133_base_resize_ack_0 : boolean;
  signal array_obj_ref_926_index_0_scale_req_0 : boolean;
  signal array_obj_ref_872_index_1_rename_req_0 : boolean;
  signal array_obj_ref_872_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_938_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_938_index_sum_1_req_1 : boolean;
  signal array_obj_ref_956_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_872_index_sum_1_req_0 : boolean;
  signal array_obj_ref_926_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_872_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_926_index_0_resize_req_0 : boolean;
  signal array_obj_ref_872_index_sum_1_req_1 : boolean;
  signal array_obj_ref_872_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_872_offset_inst_req_0 : boolean;
  signal array_obj_ref_872_offset_inst_ack_0 : boolean;
  signal array_obj_ref_950_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_938_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_944_offset_inst_ack_0 : boolean;
  signal array_obj_ref_938_index_sum_1_req_0 : boolean;
  signal array_obj_ref_872_root_address_inst_req_0 : boolean;
  signal array_obj_ref_872_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_950_index_sum_1_req_1 : boolean;
  signal array_obj_ref_944_offset_inst_req_0 : boolean;
  signal array_obj_ref_956_index_1_resize_req_0 : boolean;
  signal addr_of_873_final_reg_req_0 : boolean;
  signal addr_of_873_final_reg_ack_0 : boolean;
  signal array_obj_ref_938_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_944_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_950_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_938_index_1_rename_req_0 : boolean;
  signal array_obj_ref_944_index_sum_1_req_1 : boolean;
  signal array_obj_ref_950_index_sum_1_req_0 : boolean;
  signal array_obj_ref_944_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_938_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_938_index_1_resize_req_0 : boolean;
  signal array_obj_ref_944_index_sum_1_req_0 : boolean;
  signal binary_879_inst_req_0 : boolean;
  signal binary_879_inst_ack_0 : boolean;
  signal binary_921_inst_ack_1 : boolean;
  signal binary_879_inst_req_1 : boolean;
  signal binary_921_inst_req_1 : boolean;
  signal binary_879_inst_ack_1 : boolean;
  signal array_obj_ref_944_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_944_index_1_rename_req_0 : boolean;
  signal array_obj_ref_938_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1046_root_address_inst_req_0 : boolean;
  signal array_obj_ref_938_index_0_scale_req_1 : boolean;
  signal array_obj_ref_944_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_938_index_0_scale_ack_0 : boolean;
  signal binary_921_inst_ack_0 : boolean;
  signal binary_921_inst_req_0 : boolean;
  signal array_obj_ref_950_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_938_index_0_scale_req_0 : boolean;
  signal array_obj_ref_944_index_1_resize_req_0 : boolean;
  signal array_obj_ref_950_index_1_rename_req_0 : boolean;
  signal array_obj_ref_938_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_938_index_0_resize_req_0 : boolean;
  signal array_obj_ref_884_index_0_resize_req_0 : boolean;
  signal array_obj_ref_884_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_884_index_0_scale_req_0 : boolean;
  signal array_obj_ref_884_index_0_scale_ack_0 : boolean;
  signal addr_of_915_final_reg_ack_0 : boolean;
  signal array_obj_ref_884_index_0_scale_req_1 : boolean;
  signal addr_of_915_final_reg_req_0 : boolean;
  signal array_obj_ref_884_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1046_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_884_index_1_resize_req_0 : boolean;
  signal array_obj_ref_884_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_884_index_1_rename_req_0 : boolean;
  signal array_obj_ref_884_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_884_index_sum_1_req_0 : boolean;
  signal array_obj_ref_884_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_884_index_sum_1_req_1 : boolean;
  signal array_obj_ref_884_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_884_offset_inst_req_0 : boolean;
  signal array_obj_ref_884_offset_inst_ack_0 : boolean;
  signal array_obj_ref_884_root_address_inst_req_0 : boolean;
  signal array_obj_ref_884_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1052_root_address_inst_ack_0 : boolean;
  signal addr_of_885_final_reg_req_0 : boolean;
  signal addr_of_885_final_reg_ack_0 : boolean;
  signal array_obj_ref_1040_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1046_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1052_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1040_index_0_resize_ack_0 : boolean;
  signal addr_of_1047_final_reg_req_0 : boolean;
  signal array_obj_ref_1046_offset_inst_req_0 : boolean;
  signal array_obj_ref_1046_index_0_resize_req_0 : boolean;
  signal binary_891_inst_req_0 : boolean;
  signal array_obj_ref_1040_index_0_scale_req_0 : boolean;
  signal binary_891_inst_ack_0 : boolean;
  signal array_obj_ref_1040_index_0_scale_ack_0 : boolean;
  signal binary_891_inst_req_1 : boolean;
  signal binary_891_inst_ack_1 : boolean;
  signal array_obj_ref_1052_offset_inst_ack_0 : boolean;
  signal addr_of_1047_final_reg_ack_0 : boolean;
  signal array_obj_ref_1040_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1040_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1046_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1052_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1046_offset_inst_ack_0 : boolean;
  signal array_obj_ref_896_index_0_resize_req_0 : boolean;
  signal array_obj_ref_896_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_896_index_0_scale_req_0 : boolean;
  signal array_obj_ref_896_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_896_index_0_scale_req_1 : boolean;
  signal array_obj_ref_896_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1046_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1040_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1046_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1040_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1052_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_896_index_1_resize_req_0 : boolean;
  signal array_obj_ref_896_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_896_index_1_rename_req_0 : boolean;
  signal array_obj_ref_896_index_1_rename_ack_0 : boolean;
  signal addr_of_1053_final_reg_req_0 : boolean;
  signal array_obj_ref_1046_index_0_scale_req_1 : boolean;
  signal array_obj_ref_896_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1040_index_1_rename_req_0 : boolean;
  signal array_obj_ref_896_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_896_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1040_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_896_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_896_offset_inst_req_0 : boolean;
  signal array_obj_ref_896_offset_inst_ack_0 : boolean;
  signal addr_of_1053_final_reg_ack_0 : boolean;
  signal array_obj_ref_896_root_address_inst_req_0 : boolean;
  signal array_obj_ref_896_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1046_index_0_scale_ack_1 : boolean;
  signal addr_of_897_final_reg_req_0 : boolean;
  signal addr_of_897_final_reg_ack_0 : boolean;
  signal array_obj_ref_1052_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1052_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1052_offset_inst_req_0 : boolean;
  signal array_obj_ref_1040_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1040_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1040_index_sum_1_req_1 : boolean;
  signal array_obj_ref_902_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1040_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_902_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1052_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1040_offset_inst_req_0 : boolean;
  signal array_obj_ref_902_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1040_offset_inst_ack_0 : boolean;
  signal array_obj_ref_902_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_902_index_0_scale_req_1 : boolean;
  signal array_obj_ref_902_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_962_index_1_rename_req_0 : boolean;
  signal ptr_deref_1125_addr_0_ack_0 : boolean;
  signal array_obj_ref_962_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1052_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1040_root_address_inst_req_0 : boolean;
  signal array_obj_ref_902_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1040_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_902_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_902_index_1_rename_req_0 : boolean;
  signal array_obj_ref_902_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_902_index_sum_1_req_0 : boolean;
  signal array_obj_ref_902_index_sum_1_ack_0 : boolean;
  signal addr_of_1041_final_reg_req_0 : boolean;
  signal array_obj_ref_902_index_sum_1_req_1 : boolean;
  signal array_obj_ref_902_index_sum_1_ack_1 : boolean;
  signal addr_of_1041_final_reg_ack_0 : boolean;
  signal array_obj_ref_902_offset_inst_req_0 : boolean;
  signal array_obj_ref_902_offset_inst_ack_0 : boolean;
  signal array_obj_ref_902_root_address_inst_req_0 : boolean;
  signal array_obj_ref_902_root_address_inst_ack_0 : boolean;
  signal addr_of_903_final_reg_req_0 : boolean;
  signal addr_of_903_final_reg_ack_0 : boolean;
  signal array_obj_ref_908_index_0_resize_req_0 : boolean;
  signal array_obj_ref_908_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_908_index_0_scale_req_0 : boolean;
  signal array_obj_ref_908_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_908_index_0_scale_req_1 : boolean;
  signal array_obj_ref_908_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_908_index_1_resize_req_0 : boolean;
  signal array_obj_ref_908_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_908_index_1_rename_req_0 : boolean;
  signal array_obj_ref_908_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_908_index_sum_1_req_0 : boolean;
  signal array_obj_ref_908_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_908_index_sum_1_req_1 : boolean;
  signal array_obj_ref_908_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_908_offset_inst_req_0 : boolean;
  signal array_obj_ref_908_offset_inst_ack_0 : boolean;
  signal array_obj_ref_908_root_address_inst_req_0 : boolean;
  signal array_obj_ref_908_root_address_inst_ack_0 : boolean;
  signal addr_of_909_final_reg_req_0 : boolean;
  signal addr_of_909_final_reg_ack_0 : boolean;
  signal array_obj_ref_914_index_0_resize_req_0 : boolean;
  signal array_obj_ref_914_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_914_index_0_scale_req_0 : boolean;
  signal array_obj_ref_914_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_914_index_0_scale_req_1 : boolean;
  signal array_obj_ref_914_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_914_index_1_resize_req_0 : boolean;
  signal array_obj_ref_914_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_914_index_1_rename_req_0 : boolean;
  signal array_obj_ref_914_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_914_index_sum_1_req_0 : boolean;
  signal array_obj_ref_914_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_914_index_sum_1_req_1 : boolean;
  signal array_obj_ref_914_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_914_offset_inst_req_0 : boolean;
  signal array_obj_ref_914_offset_inst_ack_0 : boolean;
  signal array_obj_ref_914_root_address_inst_req_0 : boolean;
  signal array_obj_ref_914_root_address_inst_ack_0 : boolean;
  signal binary_1153_inst_ack_1 : boolean;
  signal array_obj_ref_962_index_sum_1_req_0 : boolean;
  signal array_obj_ref_962_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_962_index_sum_1_req_1 : boolean;
  signal array_obj_ref_962_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_962_offset_inst_req_0 : boolean;
  signal array_obj_ref_962_offset_inst_ack_0 : boolean;
  signal array_obj_ref_962_root_address_inst_req_0 : boolean;
  signal array_obj_ref_962_root_address_inst_ack_0 : boolean;
  signal binary_1158_inst_req_0 : boolean;
  signal addr_of_963_final_reg_req_0 : boolean;
  signal addr_of_963_final_reg_ack_0 : boolean;
  signal ptr_deref_1133_base_resize_req_0 : boolean;
  signal ptr_deref_1125_load_0_req_0 : boolean;
  signal binary_1138_inst_ack_0 : boolean;
  signal array_obj_ref_968_index_0_resize_req_0 : boolean;
  signal array_obj_ref_968_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1125_load_0_ack_0 : boolean;
  signal array_obj_ref_968_index_0_scale_req_0 : boolean;
  signal array_obj_ref_968_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_968_index_0_scale_req_1 : boolean;
  signal array_obj_ref_968_index_0_scale_ack_1 : boolean;
  signal ptr_deref_1133_root_address_inst_req_0 : boolean;
  signal array_obj_ref_968_index_1_resize_req_0 : boolean;
  signal array_obj_ref_968_index_1_resize_ack_0 : boolean;
  signal ptr_deref_1133_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_968_index_1_rename_req_0 : boolean;
  signal array_obj_ref_968_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_968_index_sum_1_req_0 : boolean;
  signal array_obj_ref_968_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_968_index_sum_1_req_1 : boolean;
  signal array_obj_ref_968_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_968_offset_inst_req_0 : boolean;
  signal array_obj_ref_968_offset_inst_ack_0 : boolean;
  signal binary_1153_inst_req_0 : boolean;
  signal array_obj_ref_968_root_address_inst_req_0 : boolean;
  signal array_obj_ref_968_root_address_inst_ack_0 : boolean;
  signal addr_of_969_final_reg_req_0 : boolean;
  signal addr_of_969_final_reg_ack_0 : boolean;
  signal binary_1138_inst_req_1 : boolean;
  signal ptr_deref_1125_load_0_req_1 : boolean;
  signal ptr_deref_1133_addr_0_req_0 : boolean;
  signal ptr_deref_1125_load_0_ack_1 : boolean;
  signal ptr_deref_1125_gather_scatter_req_0 : boolean;
  signal ptr_deref_1133_addr_0_ack_0 : boolean;
  signal array_obj_ref_974_index_0_resize_req_0 : boolean;
  signal array_obj_ref_974_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1125_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_974_index_0_scale_req_0 : boolean;
  signal array_obj_ref_974_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_974_index_0_scale_req_1 : boolean;
  signal array_obj_ref_974_index_0_scale_ack_1 : boolean;
  signal binary_1153_inst_ack_0 : boolean;
  signal array_obj_ref_974_index_1_resize_req_0 : boolean;
  signal array_obj_ref_974_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_974_index_1_rename_req_0 : boolean;
  signal array_obj_ref_974_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_974_index_sum_1_req_0 : boolean;
  signal array_obj_ref_974_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_974_index_sum_1_req_1 : boolean;
  signal array_obj_ref_974_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_974_offset_inst_req_0 : boolean;
  signal array_obj_ref_974_offset_inst_ack_0 : boolean;
  signal array_obj_ref_974_root_address_inst_req_0 : boolean;
  signal array_obj_ref_974_root_address_inst_ack_0 : boolean;
  signal binary_1148_inst_ack_0 : boolean;
  signal addr_of_975_final_reg_req_0 : boolean;
  signal addr_of_975_final_reg_ack_0 : boolean;
  signal binary_1138_inst_ack_1 : boolean;
  signal binary_1148_inst_ack_1 : boolean;
  signal ptr_deref_1133_load_0_req_0 : boolean;
  signal ptr_deref_1129_base_resize_req_0 : boolean;
  signal ptr_deref_1129_base_resize_ack_0 : boolean;
  signal ptr_deref_1133_load_0_ack_0 : boolean;
  signal array_obj_ref_980_index_0_resize_req_0 : boolean;
  signal array_obj_ref_980_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_980_index_0_scale_req_0 : boolean;
  signal array_obj_ref_980_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_980_index_0_scale_req_1 : boolean;
  signal array_obj_ref_980_index_0_scale_ack_1 : boolean;
  signal ptr_deref_1129_root_address_inst_req_0 : boolean;
  signal ptr_deref_1129_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_980_index_1_resize_req_0 : boolean;
  signal array_obj_ref_980_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_980_index_1_rename_req_0 : boolean;
  signal array_obj_ref_980_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_980_index_sum_1_req_0 : boolean;
  signal array_obj_ref_980_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_980_index_sum_1_req_1 : boolean;
  signal ptr_deref_1129_addr_0_req_0 : boolean;
  signal array_obj_ref_980_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_980_offset_inst_req_0 : boolean;
  signal array_obj_ref_980_offset_inst_ack_0 : boolean;
  signal ptr_deref_1129_addr_0_ack_0 : boolean;
  signal array_obj_ref_980_root_address_inst_req_0 : boolean;
  signal array_obj_ref_980_root_address_inst_ack_0 : boolean;
  signal addr_of_981_final_reg_req_0 : boolean;
  signal addr_of_981_final_reg_ack_0 : boolean;
  signal ptr_deref_1133_load_0_req_1 : boolean;
  signal binary_987_inst_req_0 : boolean;
  signal binary_987_inst_ack_0 : boolean;
  signal binary_987_inst_req_1 : boolean;
  signal binary_987_inst_ack_1 : boolean;
  signal ptr_deref_1133_load_0_ack_1 : boolean;
  signal ptr_deref_1133_gather_scatter_req_0 : boolean;
  signal ptr_deref_1129_load_0_req_0 : boolean;
  signal binary_1143_inst_req_1 : boolean;
  signal ptr_deref_1129_load_0_ack_0 : boolean;
  signal binary_993_inst_req_0 : boolean;
  signal binary_993_inst_ack_0 : boolean;
  signal binary_993_inst_req_1 : boolean;
  signal binary_993_inst_ack_1 : boolean;
  signal ptr_deref_1133_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1129_load_0_req_1 : boolean;
  signal ptr_deref_1129_load_0_ack_1 : boolean;
  signal ptr_deref_1129_gather_scatter_req_0 : boolean;
  signal array_obj_ref_998_index_0_resize_req_0 : boolean;
  signal ptr_deref_1129_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_998_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_998_index_0_scale_req_0 : boolean;
  signal array_obj_ref_998_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_998_index_0_scale_req_1 : boolean;
  signal array_obj_ref_998_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_998_index_1_resize_req_0 : boolean;
  signal array_obj_ref_998_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_998_index_1_rename_req_0 : boolean;
  signal array_obj_ref_998_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_998_index_sum_1_req_0 : boolean;
  signal array_obj_ref_998_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_998_index_sum_1_req_1 : boolean;
  signal array_obj_ref_998_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_998_offset_inst_req_0 : boolean;
  signal array_obj_ref_998_offset_inst_ack_0 : boolean;
  signal binary_1138_inst_req_0 : boolean;
  signal array_obj_ref_998_root_address_inst_req_0 : boolean;
  signal array_obj_ref_998_root_address_inst_ack_0 : boolean;
  signal addr_of_999_final_reg_req_0 : boolean;
  signal addr_of_999_final_reg_ack_0 : boolean;
  signal binary_1143_inst_req_0 : boolean;
  signal binary_1158_inst_ack_0 : boolean;
  signal binary_1158_inst_req_1 : boolean;
  signal binary_1158_inst_ack_1 : boolean;
  signal binary_1005_inst_req_0 : boolean;
  signal binary_1005_inst_ack_0 : boolean;
  signal binary_1153_inst_req_1 : boolean;
  signal binary_1005_inst_req_1 : boolean;
  signal binary_1005_inst_ack_1 : boolean;
  signal binary_1143_inst_ack_0 : boolean;
  signal binary_1148_inst_req_1 : boolean;
  signal array_obj_ref_1010_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1010_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1010_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1010_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1010_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1010_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1010_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1010_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1010_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1010_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1010_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1010_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1010_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1010_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1010_offset_inst_req_0 : boolean;
  signal array_obj_ref_1010_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1010_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1010_root_address_inst_ack_0 : boolean;
  signal addr_of_1011_final_reg_req_0 : boolean;
  signal addr_of_1011_final_reg_ack_0 : boolean;
  signal binary_1017_inst_req_0 : boolean;
  signal binary_1017_inst_ack_0 : boolean;
  signal binary_1017_inst_req_1 : boolean;
  signal binary_1017_inst_ack_1 : boolean;
  signal array_obj_ref_1022_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1022_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1022_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1022_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1022_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1022_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1022_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1022_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1022_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1022_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1022_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1022_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1022_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1022_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1022_offset_inst_req_0 : boolean;
  signal array_obj_ref_1022_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1022_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1022_root_address_inst_ack_0 : boolean;
  signal addr_of_1023_final_reg_req_0 : boolean;
  signal addr_of_1023_final_reg_ack_0 : boolean;
  signal array_obj_ref_1028_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1028_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1028_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1028_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1028_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1028_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1028_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1028_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1028_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1028_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1028_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1028_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1028_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1028_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1028_offset_inst_req_0 : boolean;
  signal array_obj_ref_1028_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1028_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1028_root_address_inst_ack_0 : boolean;
  signal addr_of_1029_final_reg_req_0 : boolean;
  signal addr_of_1029_final_reg_ack_0 : boolean;
  signal array_obj_ref_1034_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1034_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1034_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1034_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1034_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1034_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1034_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1034_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1034_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1034_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1034_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1034_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1034_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1034_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1034_offset_inst_req_0 : boolean;
  signal array_obj_ref_1034_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1034_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1034_root_address_inst_ack_0 : boolean;
  signal addr_of_1035_final_reg_req_0 : boolean;
  signal addr_of_1035_final_reg_ack_0 : boolean;
  signal array_obj_ref_1058_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1058_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1058_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1058_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1058_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1058_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1058_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1058_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1058_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1058_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1058_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1058_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1058_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1058_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1058_offset_inst_req_0 : boolean;
  signal array_obj_ref_1058_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1058_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1058_root_address_inst_ack_0 : boolean;
  signal addr_of_1059_final_reg_req_0 : boolean;
  signal addr_of_1059_final_reg_ack_0 : boolean;
  signal array_obj_ref_1064_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1064_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1064_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1064_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1064_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1064_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1064_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1064_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1064_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1064_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1064_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1064_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1064_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1064_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1064_offset_inst_req_0 : boolean;
  signal array_obj_ref_1064_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1064_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1064_root_address_inst_ack_0 : boolean;
  signal addr_of_1065_final_reg_req_0 : boolean;
  signal addr_of_1065_final_reg_ack_0 : boolean;
  signal array_obj_ref_1070_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1070_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1070_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1070_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1070_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1070_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1070_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1070_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1070_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1070_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1070_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1070_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1070_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1070_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1070_offset_inst_req_0 : boolean;
  signal array_obj_ref_1070_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1070_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1070_root_address_inst_ack_0 : boolean;
  signal addr_of_1071_final_reg_req_0 : boolean;
  signal addr_of_1071_final_reg_ack_0 : boolean;
  signal binary_1280_inst_req_0 : boolean;
  signal binary_1280_inst_ack_0 : boolean;
  signal array_obj_ref_1076_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1076_index_0_resize_ack_0 : boolean;
  signal binary_1285_inst_ack_0 : boolean;
  signal array_obj_ref_1076_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1076_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1076_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1076_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1076_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1076_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1076_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1076_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1076_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1076_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1076_index_sum_1_req_1 : boolean;
  signal binary_1265_inst_req_0 : boolean;
  signal array_obj_ref_1076_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1076_offset_inst_req_0 : boolean;
  signal array_obj_ref_1076_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1076_root_address_inst_req_0 : boolean;
  signal binary_1265_inst_ack_0 : boolean;
  signal array_obj_ref_1076_root_address_inst_ack_0 : boolean;
  signal addr_of_1077_final_reg_req_0 : boolean;
  signal binary_1265_inst_req_1 : boolean;
  signal addr_of_1077_final_reg_ack_0 : boolean;
  signal binary_1265_inst_ack_1 : boolean;
  signal binary_1280_inst_req_1 : boolean;
  signal binary_1280_inst_ack_1 : boolean;
  signal binary_1285_inst_req_1 : boolean;
  signal array_obj_ref_1082_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1082_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1289_load_0_ack_1 : boolean;
  signal array_obj_ref_1082_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1082_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1082_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1082_index_0_scale_ack_1 : boolean;
  signal binary_1285_inst_ack_1 : boolean;
  signal array_obj_ref_1082_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1082_index_1_resize_ack_0 : boolean;
  signal ptr_deref_1289_addr_0_req_0 : boolean;
  signal array_obj_ref_1082_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1082_index_1_rename_ack_0 : boolean;
  signal ptr_deref_1289_load_0_req_1 : boolean;
  signal array_obj_ref_1082_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1082_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1082_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1082_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1082_offset_inst_req_0 : boolean;
  signal array_obj_ref_1082_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1082_root_address_inst_req_0 : boolean;
  signal binary_1270_inst_req_0 : boolean;
  signal array_obj_ref_1082_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1289_gather_scatter_req_0 : boolean;
  signal binary_1270_inst_ack_0 : boolean;
  signal addr_of_1083_final_reg_req_0 : boolean;
  signal addr_of_1083_final_reg_ack_0 : boolean;
  signal binary_1270_inst_req_1 : boolean;
  signal binary_1270_inst_ack_1 : boolean;
  signal ptr_deref_1289_root_address_inst_req_0 : boolean;
  signal ptr_deref_1289_load_0_req_0 : boolean;
  signal array_obj_ref_1088_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1088_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1088_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1088_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1088_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1088_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1088_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1088_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1088_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1088_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1088_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1088_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1088_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1088_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1088_offset_inst_req_0 : boolean;
  signal array_obj_ref_1088_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1088_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1088_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1289_load_0_ack_0 : boolean;
  signal addr_of_1089_final_reg_req_0 : boolean;
  signal addr_of_1089_final_reg_ack_0 : boolean;
  signal binary_1275_inst_req_0 : boolean;
  signal binary_1275_inst_ack_0 : boolean;
  signal binary_1275_inst_req_1 : boolean;
  signal ptr_deref_1289_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1094_index_0_resize_req_0 : boolean;
  signal binary_1275_inst_ack_1 : boolean;
  signal array_obj_ref_1094_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1094_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1094_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1094_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1094_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1094_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1094_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1094_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1094_index_1_rename_ack_0 : boolean;
  signal ptr_deref_1289_addr_0_ack_0 : boolean;
  signal array_obj_ref_1094_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1094_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1094_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1094_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1094_offset_inst_req_0 : boolean;
  signal array_obj_ref_1094_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1094_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1094_root_address_inst_ack_0 : boolean;
  signal addr_of_1095_final_reg_req_0 : boolean;
  signal addr_of_1095_final_reg_ack_0 : boolean;
  signal binary_1658_inst_ack_0 : boolean;
  signal binary_1285_inst_req_0 : boolean;
  signal ptr_deref_1289_base_resize_req_0 : boolean;
  signal array_obj_ref_1100_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1100_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1100_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1100_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1100_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1100_index_0_scale_ack_1 : boolean;
  signal ptr_deref_1289_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1289_base_resize_ack_0 : boolean;
  signal array_obj_ref_1100_index_1_resize_req_0 : boolean;
  signal array_obj_ref_1100_index_1_resize_ack_0 : boolean;
  signal array_obj_ref_1100_index_1_rename_req_0 : boolean;
  signal array_obj_ref_1100_index_1_rename_ack_0 : boolean;
  signal array_obj_ref_1100_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1100_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1100_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1100_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1100_offset_inst_req_0 : boolean;
  signal array_obj_ref_1100_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1100_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1100_root_address_inst_ack_0 : boolean;
  signal addr_of_1101_final_reg_req_0 : boolean;
  signal addr_of_1101_final_reg_ack_0 : boolean;
  signal ptr_deref_1105_base_resize_req_0 : boolean;
  signal ptr_deref_1105_base_resize_ack_0 : boolean;
  signal ptr_deref_1105_root_address_inst_req_0 : boolean;
  signal ptr_deref_1105_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1105_addr_0_req_0 : boolean;
  signal ptr_deref_1105_addr_0_ack_0 : boolean;
  signal ptr_deref_1105_load_0_req_0 : boolean;
  signal ptr_deref_1105_load_0_ack_0 : boolean;
  signal ptr_deref_1105_load_0_req_1 : boolean;
  signal ptr_deref_1105_load_0_ack_1 : boolean;
  signal ptr_deref_1105_gather_scatter_req_0 : boolean;
  signal ptr_deref_1105_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1109_base_resize_req_0 : boolean;
  signal ptr_deref_1109_base_resize_ack_0 : boolean;
  signal ptr_deref_1109_root_address_inst_req_0 : boolean;
  signal ptr_deref_1109_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1109_addr_0_req_0 : boolean;
  signal ptr_deref_1109_addr_0_ack_0 : boolean;
  signal ptr_deref_1109_load_0_req_0 : boolean;
  signal ptr_deref_1109_load_0_ack_0 : boolean;
  signal ptr_deref_1109_load_0_req_1 : boolean;
  signal ptr_deref_1109_load_0_ack_1 : boolean;
  signal ptr_deref_1109_gather_scatter_req_0 : boolean;
  signal ptr_deref_1109_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1113_base_resize_req_0 : boolean;
  signal ptr_deref_1113_base_resize_ack_0 : boolean;
  signal ptr_deref_1113_root_address_inst_req_0 : boolean;
  signal ptr_deref_1113_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1113_addr_0_req_0 : boolean;
  signal ptr_deref_1113_addr_0_ack_0 : boolean;
  signal ptr_deref_1113_load_0_req_0 : boolean;
  signal ptr_deref_1113_load_0_ack_0 : boolean;
  signal ptr_deref_1113_load_0_req_1 : boolean;
  signal ptr_deref_1113_load_0_ack_1 : boolean;
  signal ptr_deref_1113_gather_scatter_req_0 : boolean;
  signal ptr_deref_1113_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1117_base_resize_req_0 : boolean;
  signal ptr_deref_1117_base_resize_ack_0 : boolean;
  signal ptr_deref_1117_root_address_inst_req_0 : boolean;
  signal ptr_deref_1117_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1117_addr_0_req_0 : boolean;
  signal ptr_deref_1117_addr_0_ack_0 : boolean;
  signal ptr_deref_1117_load_0_req_0 : boolean;
  signal ptr_deref_1117_load_0_ack_0 : boolean;
  signal ptr_deref_1117_load_0_req_1 : boolean;
  signal ptr_deref_1117_load_0_ack_1 : boolean;
  signal ptr_deref_1117_gather_scatter_req_0 : boolean;
  signal ptr_deref_1117_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1121_base_resize_req_0 : boolean;
  signal ptr_deref_1121_base_resize_ack_0 : boolean;
  signal ptr_deref_1121_root_address_inst_req_0 : boolean;
  signal ptr_deref_1121_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1121_addr_0_req_0 : boolean;
  signal ptr_deref_1121_addr_0_ack_0 : boolean;
  signal ptr_deref_1121_load_0_req_0 : boolean;
  signal ptr_deref_1121_load_0_ack_0 : boolean;
  signal ptr_deref_1121_load_0_req_1 : boolean;
  signal ptr_deref_1121_load_0_ack_1 : boolean;
  signal ptr_deref_1121_gather_scatter_req_0 : boolean;
  signal ptr_deref_1121_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1125_base_resize_req_0 : boolean;
  signal ptr_deref_1125_base_resize_ack_0 : boolean;
  signal ptr_deref_1125_root_address_inst_req_0 : boolean;
  signal ptr_deref_1125_root_address_inst_ack_0 : boolean;
  signal binary_1447_inst_req_0 : boolean;
  signal binary_1447_inst_ack_0 : boolean;
  signal binary_1447_inst_req_1 : boolean;
  signal binary_1447_inst_ack_1 : boolean;
  signal binary_1163_inst_req_0 : boolean;
  signal binary_1163_inst_ack_0 : boolean;
  signal binary_1163_inst_req_1 : boolean;
  signal binary_1163_inst_ack_1 : boolean;
  signal binary_1168_inst_req_0 : boolean;
  signal binary_1168_inst_ack_0 : boolean;
  signal binary_1168_inst_req_1 : boolean;
  signal binary_1168_inst_ack_1 : boolean;
  signal binary_1173_inst_req_0 : boolean;
  signal binary_1173_inst_ack_0 : boolean;
  signal binary_1173_inst_req_1 : boolean;
  signal binary_1173_inst_ack_1 : boolean;
  signal ptr_deref_1177_base_resize_req_0 : boolean;
  signal ptr_deref_1177_base_resize_ack_0 : boolean;
  signal ptr_deref_1177_root_address_inst_req_0 : boolean;
  signal ptr_deref_1177_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1177_addr_0_req_0 : boolean;
  signal ptr_deref_1177_addr_0_ack_0 : boolean;
  signal ptr_deref_1177_load_0_req_0 : boolean;
  signal ptr_deref_1177_load_0_ack_0 : boolean;
  signal ptr_deref_1177_load_0_req_1 : boolean;
  signal ptr_deref_1177_load_0_ack_1 : boolean;
  signal ptr_deref_1177_gather_scatter_req_0 : boolean;
  signal ptr_deref_1177_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1181_base_resize_req_0 : boolean;
  signal ptr_deref_1181_base_resize_ack_0 : boolean;
  signal ptr_deref_1181_root_address_inst_req_0 : boolean;
  signal ptr_deref_1181_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1181_addr_0_req_0 : boolean;
  signal ptr_deref_1181_addr_0_ack_0 : boolean;
  signal ptr_deref_1181_load_0_req_0 : boolean;
  signal ptr_deref_1181_load_0_ack_0 : boolean;
  signal ptr_deref_1181_load_0_req_1 : boolean;
  signal ptr_deref_1181_load_0_ack_1 : boolean;
  signal ptr_deref_1181_gather_scatter_req_0 : boolean;
  signal ptr_deref_1181_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1185_base_resize_req_0 : boolean;
  signal ptr_deref_1185_base_resize_ack_0 : boolean;
  signal ptr_deref_1185_root_address_inst_req_0 : boolean;
  signal ptr_deref_1185_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1185_addr_0_req_0 : boolean;
  signal ptr_deref_1185_addr_0_ack_0 : boolean;
  signal ptr_deref_1185_load_0_req_0 : boolean;
  signal ptr_deref_1185_load_0_ack_0 : boolean;
  signal ptr_deref_1185_load_0_req_1 : boolean;
  signal ptr_deref_1185_load_0_ack_1 : boolean;
  signal ptr_deref_1185_gather_scatter_req_0 : boolean;
  signal ptr_deref_1185_gather_scatter_ack_0 : boolean;
  signal binary_1643_inst_req_0 : boolean;
  signal ptr_deref_1189_base_resize_req_0 : boolean;
  signal ptr_deref_1189_base_resize_ack_0 : boolean;
  signal ptr_deref_1189_root_address_inst_req_0 : boolean;
  signal ptr_deref_1189_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1189_addr_0_req_0 : boolean;
  signal ptr_deref_1189_addr_0_ack_0 : boolean;
  signal ptr_deref_1189_load_0_req_0 : boolean;
  signal ptr_deref_1189_load_0_ack_0 : boolean;
  signal binary_1633_inst_req_1 : boolean;
  signal ptr_deref_1189_load_0_req_1 : boolean;
  signal ptr_deref_1189_load_0_ack_1 : boolean;
  signal ptr_deref_1189_gather_scatter_req_0 : boolean;
  signal ptr_deref_1189_gather_scatter_ack_0 : boolean;
  signal binary_1643_inst_ack_0 : boolean;
  signal binary_1194_inst_req_0 : boolean;
  signal binary_1194_inst_ack_0 : boolean;
  signal binary_1194_inst_req_1 : boolean;
  signal binary_1194_inst_ack_1 : boolean;
  signal binary_1407_inst_req_0 : boolean;
  signal binary_1407_inst_ack_0 : boolean;
  signal binary_1633_inst_ack_1 : boolean;
  signal binary_1199_inst_req_0 : boolean;
  signal binary_1199_inst_ack_0 : boolean;
  signal binary_1199_inst_req_1 : boolean;
  signal binary_1199_inst_ack_1 : boolean;
  signal binary_1204_inst_req_0 : boolean;
  signal binary_1204_inst_ack_0 : boolean;
  signal binary_1204_inst_req_1 : boolean;
  signal binary_1204_inst_ack_1 : boolean;
  signal binary_1209_inst_req_0 : boolean;
  signal binary_1209_inst_ack_0 : boolean;
  signal binary_1209_inst_req_1 : boolean;
  signal binary_1209_inst_ack_1 : boolean;
  signal binary_1214_inst_req_0 : boolean;
  signal binary_1214_inst_ack_0 : boolean;
  signal binary_1214_inst_req_1 : boolean;
  signal binary_1214_inst_ack_1 : boolean;
  signal binary_1219_inst_req_0 : boolean;
  signal binary_1219_inst_ack_0 : boolean;
  signal binary_1219_inst_req_1 : boolean;
  signal binary_1219_inst_ack_1 : boolean;
  signal binary_1224_inst_req_0 : boolean;
  signal binary_1224_inst_ack_0 : boolean;
  signal binary_1224_inst_req_1 : boolean;
  signal binary_1224_inst_ack_1 : boolean;
  signal binary_1229_inst_req_0 : boolean;
  signal binary_1229_inst_ack_0 : boolean;
  signal binary_1229_inst_req_1 : boolean;
  signal binary_1229_inst_ack_1 : boolean;
  signal ptr_deref_1233_base_resize_req_0 : boolean;
  signal ptr_deref_1233_base_resize_ack_0 : boolean;
  signal ptr_deref_1233_root_address_inst_req_0 : boolean;
  signal ptr_deref_1233_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1233_addr_0_req_0 : boolean;
  signal ptr_deref_1233_addr_0_ack_0 : boolean;
  signal ptr_deref_1233_load_0_req_0 : boolean;
  signal ptr_deref_1233_load_0_ack_0 : boolean;
  signal ptr_deref_1233_load_0_req_1 : boolean;
  signal ptr_deref_1233_load_0_ack_1 : boolean;
  signal ptr_deref_1233_gather_scatter_req_0 : boolean;
  signal ptr_deref_1233_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1237_base_resize_req_0 : boolean;
  signal ptr_deref_1237_base_resize_ack_0 : boolean;
  signal ptr_deref_1237_root_address_inst_req_0 : boolean;
  signal ptr_deref_1237_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1237_addr_0_req_0 : boolean;
  signal ptr_deref_1237_addr_0_ack_0 : boolean;
  signal ptr_deref_1237_load_0_req_0 : boolean;
  signal ptr_deref_1237_load_0_ack_0 : boolean;
  signal ptr_deref_1237_load_0_req_1 : boolean;
  signal ptr_deref_1237_load_0_ack_1 : boolean;
  signal ptr_deref_1237_gather_scatter_req_0 : boolean;
  signal ptr_deref_1237_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1241_base_resize_req_0 : boolean;
  signal ptr_deref_1241_base_resize_ack_0 : boolean;
  signal ptr_deref_1241_root_address_inst_req_0 : boolean;
  signal ptr_deref_1241_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1241_addr_0_req_0 : boolean;
  signal ptr_deref_1241_addr_0_ack_0 : boolean;
  signal ptr_deref_1241_load_0_req_0 : boolean;
  signal ptr_deref_1241_load_0_ack_0 : boolean;
  signal ptr_deref_1241_load_0_req_1 : boolean;
  signal ptr_deref_1241_load_0_ack_1 : boolean;
  signal ptr_deref_1241_gather_scatter_req_0 : boolean;
  signal ptr_deref_1241_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1245_base_resize_req_0 : boolean;
  signal ptr_deref_1245_base_resize_ack_0 : boolean;
  signal ptr_deref_1245_root_address_inst_req_0 : boolean;
  signal ptr_deref_1245_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1245_addr_0_req_0 : boolean;
  signal ptr_deref_1245_addr_0_ack_0 : boolean;
  signal ptr_deref_1245_load_0_req_0 : boolean;
  signal ptr_deref_1245_load_0_ack_0 : boolean;
  signal ptr_deref_1245_load_0_req_1 : boolean;
  signal ptr_deref_1245_load_0_ack_1 : boolean;
  signal ptr_deref_1245_gather_scatter_req_0 : boolean;
  signal ptr_deref_1245_gather_scatter_ack_0 : boolean;
  signal binary_1250_inst_req_0 : boolean;
  signal binary_1250_inst_ack_0 : boolean;
  signal binary_1250_inst_req_1 : boolean;
  signal binary_1250_inst_ack_1 : boolean;
  signal binary_1255_inst_req_0 : boolean;
  signal binary_1255_inst_ack_0 : boolean;
  signal binary_1255_inst_req_1 : boolean;
  signal binary_1255_inst_ack_1 : boolean;
  signal binary_1260_inst_req_0 : boolean;
  signal binary_1260_inst_ack_0 : boolean;
  signal binary_1260_inst_req_1 : boolean;
  signal binary_1260_inst_ack_1 : boolean;
  signal ptr_deref_1293_base_resize_req_0 : boolean;
  signal ptr_deref_1293_base_resize_ack_0 : boolean;
  signal ptr_deref_1293_root_address_inst_req_0 : boolean;
  signal ptr_deref_1293_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1293_addr_0_req_0 : boolean;
  signal ptr_deref_1293_addr_0_ack_0 : boolean;
  signal ptr_deref_1293_load_0_req_0 : boolean;
  signal ptr_deref_1293_load_0_ack_0 : boolean;
  signal ptr_deref_1293_load_0_req_1 : boolean;
  signal ptr_deref_1293_load_0_ack_1 : boolean;
  signal ptr_deref_1293_gather_scatter_req_0 : boolean;
  signal ptr_deref_1293_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1297_base_resize_req_0 : boolean;
  signal ptr_deref_1297_base_resize_ack_0 : boolean;
  signal ptr_deref_1297_root_address_inst_req_0 : boolean;
  signal ptr_deref_1297_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1297_addr_0_req_0 : boolean;
  signal ptr_deref_1297_addr_0_ack_0 : boolean;
  signal ptr_deref_1297_load_0_req_0 : boolean;
  signal ptr_deref_1297_load_0_ack_0 : boolean;
  signal ptr_deref_1297_load_0_req_1 : boolean;
  signal ptr_deref_1297_load_0_ack_1 : boolean;
  signal ptr_deref_1297_gather_scatter_req_0 : boolean;
  signal ptr_deref_1297_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1301_base_resize_req_0 : boolean;
  signal ptr_deref_1301_base_resize_ack_0 : boolean;
  signal ptr_deref_1301_root_address_inst_req_0 : boolean;
  signal ptr_deref_1301_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1301_addr_0_req_0 : boolean;
  signal ptr_deref_1301_addr_0_ack_0 : boolean;
  signal ptr_deref_1301_load_0_req_0 : boolean;
  signal ptr_deref_1301_load_0_ack_0 : boolean;
  signal ptr_deref_1301_load_0_req_1 : boolean;
  signal ptr_deref_1301_load_0_ack_1 : boolean;
  signal ptr_deref_1301_gather_scatter_req_0 : boolean;
  signal ptr_deref_1301_gather_scatter_ack_0 : boolean;
  signal binary_1306_inst_req_0 : boolean;
  signal binary_1306_inst_ack_0 : boolean;
  signal binary_1306_inst_req_1 : boolean;
  signal binary_1306_inst_ack_1 : boolean;
  signal binary_1311_inst_req_0 : boolean;
  signal binary_1311_inst_ack_0 : boolean;
  signal binary_1311_inst_req_1 : boolean;
  signal binary_1311_inst_ack_1 : boolean;
  signal binary_1316_inst_req_0 : boolean;
  signal binary_1316_inst_ack_0 : boolean;
  signal binary_1316_inst_req_1 : boolean;
  signal binary_1316_inst_ack_1 : boolean;
  signal binary_1321_inst_req_0 : boolean;
  signal binary_1321_inst_ack_0 : boolean;
  signal binary_1321_inst_req_1 : boolean;
  signal binary_1321_inst_ack_1 : boolean;
  signal binary_1326_inst_req_0 : boolean;
  signal binary_1326_inst_ack_0 : boolean;
  signal binary_1326_inst_req_1 : boolean;
  signal binary_1326_inst_ack_1 : boolean;
  signal binary_1331_inst_req_0 : boolean;
  signal binary_1331_inst_ack_0 : boolean;
  signal binary_1331_inst_req_1 : boolean;
  signal binary_1331_inst_ack_1 : boolean;
  signal binary_1336_inst_req_0 : boolean;
  signal binary_1336_inst_ack_0 : boolean;
  signal binary_1336_inst_req_1 : boolean;
  signal binary_1336_inst_ack_1 : boolean;
  signal binary_1341_inst_req_0 : boolean;
  signal binary_1341_inst_ack_0 : boolean;
  signal binary_1341_inst_req_1 : boolean;
  signal binary_1341_inst_ack_1 : boolean;
  signal ptr_deref_1345_base_resize_req_0 : boolean;
  signal ptr_deref_1345_base_resize_ack_0 : boolean;
  signal ptr_deref_1345_root_address_inst_req_0 : boolean;
  signal ptr_deref_1345_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1345_addr_0_req_0 : boolean;
  signal ptr_deref_1345_addr_0_ack_0 : boolean;
  signal ptr_deref_1345_load_0_req_0 : boolean;
  signal ptr_deref_1345_load_0_ack_0 : boolean;
  signal ptr_deref_1345_load_0_req_1 : boolean;
  signal ptr_deref_1345_load_0_ack_1 : boolean;
  signal ptr_deref_1345_gather_scatter_req_0 : boolean;
  signal ptr_deref_1345_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1349_base_resize_req_0 : boolean;
  signal ptr_deref_1349_base_resize_ack_0 : boolean;
  signal ptr_deref_1349_root_address_inst_req_0 : boolean;
  signal ptr_deref_1349_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1349_addr_0_req_0 : boolean;
  signal ptr_deref_1349_addr_0_ack_0 : boolean;
  signal ptr_deref_1349_load_0_req_0 : boolean;
  signal ptr_deref_1349_load_0_ack_0 : boolean;
  signal ptr_deref_1349_load_0_req_1 : boolean;
  signal ptr_deref_1349_load_0_ack_1 : boolean;
  signal ptr_deref_1349_gather_scatter_req_0 : boolean;
  signal ptr_deref_1349_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1353_base_resize_req_0 : boolean;
  signal ptr_deref_1353_base_resize_ack_0 : boolean;
  signal ptr_deref_1353_root_address_inst_req_0 : boolean;
  signal ptr_deref_1353_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1353_addr_0_req_0 : boolean;
  signal ptr_deref_1353_addr_0_ack_0 : boolean;
  signal ptr_deref_1353_load_0_req_0 : boolean;
  signal ptr_deref_1353_load_0_ack_0 : boolean;
  signal ptr_deref_1353_load_0_req_1 : boolean;
  signal ptr_deref_1353_load_0_ack_1 : boolean;
  signal ptr_deref_1353_gather_scatter_req_0 : boolean;
  signal ptr_deref_1353_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1357_base_resize_req_0 : boolean;
  signal ptr_deref_1357_base_resize_ack_0 : boolean;
  signal ptr_deref_1357_root_address_inst_req_0 : boolean;
  signal ptr_deref_1357_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1357_addr_0_req_0 : boolean;
  signal ptr_deref_1357_addr_0_ack_0 : boolean;
  signal ptr_deref_1357_load_0_req_0 : boolean;
  signal ptr_deref_1357_load_0_ack_0 : boolean;
  signal ptr_deref_1357_load_0_req_1 : boolean;
  signal ptr_deref_1357_load_0_ack_1 : boolean;
  signal ptr_deref_1357_gather_scatter_req_0 : boolean;
  signal ptr_deref_1357_gather_scatter_ack_0 : boolean;
  signal binary_1362_inst_req_0 : boolean;
  signal binary_1362_inst_ack_0 : boolean;
  signal binary_1362_inst_req_1 : boolean;
  signal binary_1362_inst_ack_1 : boolean;
  signal binary_1367_inst_req_0 : boolean;
  signal binary_1367_inst_ack_0 : boolean;
  signal binary_1367_inst_req_1 : boolean;
  signal binary_1367_inst_ack_1 : boolean;
  signal binary_1372_inst_req_0 : boolean;
  signal binary_1372_inst_ack_0 : boolean;
  signal binary_1372_inst_req_1 : boolean;
  signal binary_1372_inst_ack_1 : boolean;
  signal binary_1377_inst_req_0 : boolean;
  signal binary_1377_inst_ack_0 : boolean;
  signal binary_1377_inst_req_1 : boolean;
  signal binary_1377_inst_ack_1 : boolean;
  signal binary_1382_inst_req_0 : boolean;
  signal binary_1382_inst_ack_0 : boolean;
  signal binary_1382_inst_req_1 : boolean;
  signal binary_1382_inst_ack_1 : boolean;
  signal binary_1387_inst_req_0 : boolean;
  signal binary_1387_inst_ack_0 : boolean;
  signal binary_1387_inst_req_1 : boolean;
  signal binary_1387_inst_ack_1 : boolean;
  signal binary_1392_inst_req_0 : boolean;
  signal binary_1392_inst_ack_0 : boolean;
  signal binary_1392_inst_req_1 : boolean;
  signal binary_1392_inst_ack_1 : boolean;
  signal binary_1397_inst_req_0 : boolean;
  signal binary_1397_inst_ack_0 : boolean;
  signal binary_1397_inst_req_1 : boolean;
  signal binary_1397_inst_ack_1 : boolean;
  signal binary_1402_inst_req_0 : boolean;
  signal binary_1402_inst_ack_0 : boolean;
  signal binary_1402_inst_req_1 : boolean;
  signal binary_1402_inst_ack_1 : boolean;
  signal binary_1407_inst_req_1 : boolean;
  signal binary_1407_inst_ack_1 : boolean;
  signal binary_1412_inst_req_0 : boolean;
  signal binary_1412_inst_ack_0 : boolean;
  signal binary_1412_inst_req_1 : boolean;
  signal binary_1412_inst_ack_1 : boolean;
  signal binary_1417_inst_req_0 : boolean;
  signal binary_1417_inst_ack_0 : boolean;
  signal binary_1417_inst_req_1 : boolean;
  signal binary_1417_inst_ack_1 : boolean;
  signal binary_1422_inst_req_0 : boolean;
  signal binary_1422_inst_ack_0 : boolean;
  signal binary_1422_inst_req_1 : boolean;
  signal binary_1422_inst_ack_1 : boolean;
  signal binary_1663_inst_ack_0 : boolean;
  signal binary_1643_inst_req_1 : boolean;
  signal binary_1653_inst_req_0 : boolean;
  signal binary_1427_inst_req_0 : boolean;
  signal binary_1427_inst_ack_0 : boolean;
  signal binary_1427_inst_req_1 : boolean;
  signal binary_1427_inst_ack_1 : boolean;
  signal binary_1643_inst_ack_1 : boolean;
  signal binary_1658_inst_req_1 : boolean;
  signal binary_1653_inst_req_1 : boolean;
  signal binary_1653_inst_ack_1 : boolean;
  signal binary_1638_inst_req_0 : boolean;
  signal binary_1432_inst_req_0 : boolean;
  signal binary_1432_inst_ack_0 : boolean;
  signal binary_1432_inst_req_1 : boolean;
  signal binary_1432_inst_ack_1 : boolean;
  signal binary_1638_inst_ack_0 : boolean;
  signal binary_1663_inst_req_0 : boolean;
  signal binary_1638_inst_req_1 : boolean;
  signal binary_1658_inst_req_0 : boolean;
  signal binary_1638_inst_ack_1 : boolean;
  signal binary_1437_inst_req_0 : boolean;
  signal binary_1437_inst_ack_0 : boolean;
  signal binary_1437_inst_req_1 : boolean;
  signal binary_1437_inst_ack_1 : boolean;
  signal binary_1663_inst_req_1 : boolean;
  signal binary_1442_inst_req_0 : boolean;
  signal binary_1442_inst_ack_0 : boolean;
  signal binary_1442_inst_req_1 : boolean;
  signal binary_1442_inst_ack_1 : boolean;
  signal binary_1648_inst_req_0 : boolean;
  signal binary_1648_inst_ack_0 : boolean;
  signal binary_1653_inst_ack_0 : boolean;
  signal binary_1648_inst_req_1 : boolean;
  signal binary_1658_inst_ack_1 : boolean;
  signal binary_1648_inst_ack_1 : boolean;
  signal binary_1452_inst_req_0 : boolean;
  signal binary_1452_inst_ack_0 : boolean;
  signal binary_1452_inst_req_1 : boolean;
  signal binary_1452_inst_ack_1 : boolean;
  signal binary_1663_inst_ack_1 : boolean;
  signal binary_1457_inst_req_0 : boolean;
  signal binary_1457_inst_ack_0 : boolean;
  signal binary_1457_inst_req_1 : boolean;
  signal binary_1457_inst_ack_1 : boolean;
  signal binary_1462_inst_req_0 : boolean;
  signal binary_1462_inst_ack_0 : boolean;
  signal binary_1462_inst_req_1 : boolean;
  signal binary_1462_inst_ack_1 : boolean;
  signal binary_1467_inst_req_0 : boolean;
  signal binary_1467_inst_ack_0 : boolean;
  signal binary_1467_inst_req_1 : boolean;
  signal binary_1467_inst_ack_1 : boolean;
  signal binary_1472_inst_req_0 : boolean;
  signal binary_1472_inst_ack_0 : boolean;
  signal binary_1472_inst_req_1 : boolean;
  signal binary_1472_inst_ack_1 : boolean;
  signal binary_1477_inst_req_0 : boolean;
  signal binary_1477_inst_ack_0 : boolean;
  signal binary_1477_inst_req_1 : boolean;
  signal binary_1477_inst_ack_1 : boolean;
  signal binary_1482_inst_req_0 : boolean;
  signal binary_1482_inst_ack_0 : boolean;
  signal binary_1482_inst_req_1 : boolean;
  signal binary_1482_inst_ack_1 : boolean;
  signal binary_1487_inst_req_0 : boolean;
  signal binary_1487_inst_ack_0 : boolean;
  signal binary_1487_inst_req_1 : boolean;
  signal binary_1487_inst_ack_1 : boolean;
  signal binary_1492_inst_req_0 : boolean;
  signal binary_1492_inst_ack_0 : boolean;
  signal binary_1492_inst_req_1 : boolean;
  signal binary_1492_inst_ack_1 : boolean;
  signal binary_1497_inst_req_0 : boolean;
  signal binary_1497_inst_ack_0 : boolean;
  signal binary_1497_inst_req_1 : boolean;
  signal binary_1497_inst_ack_1 : boolean;
  signal binary_1502_inst_req_0 : boolean;
  signal binary_1502_inst_ack_0 : boolean;
  signal binary_1502_inst_req_1 : boolean;
  signal binary_1502_inst_ack_1 : boolean;
  signal binary_1507_inst_req_0 : boolean;
  signal binary_1507_inst_ack_0 : boolean;
  signal binary_1507_inst_req_1 : boolean;
  signal binary_1507_inst_ack_1 : boolean;
  signal binary_1512_inst_req_0 : boolean;
  signal binary_1512_inst_ack_0 : boolean;
  signal binary_1512_inst_req_1 : boolean;
  signal binary_1512_inst_ack_1 : boolean;
  signal binary_1517_inst_req_0 : boolean;
  signal binary_1517_inst_ack_0 : boolean;
  signal binary_1517_inst_req_1 : boolean;
  signal binary_1517_inst_ack_1 : boolean;
  signal ptr_deref_1521_base_resize_req_0 : boolean;
  signal ptr_deref_1521_base_resize_ack_0 : boolean;
  signal ptr_deref_1521_root_address_inst_req_0 : boolean;
  signal ptr_deref_1521_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1521_addr_0_req_0 : boolean;
  signal ptr_deref_1521_addr_0_ack_0 : boolean;
  signal ptr_deref_1521_load_0_req_0 : boolean;
  signal ptr_deref_1521_load_0_ack_0 : boolean;
  signal ptr_deref_1521_load_0_req_1 : boolean;
  signal ptr_deref_1521_load_0_ack_1 : boolean;
  signal ptr_deref_1521_gather_scatter_req_0 : boolean;
  signal ptr_deref_1521_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1525_base_resize_req_0 : boolean;
  signal ptr_deref_1525_base_resize_ack_0 : boolean;
  signal ptr_deref_1525_root_address_inst_req_0 : boolean;
  signal ptr_deref_1525_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1525_addr_0_req_0 : boolean;
  signal ptr_deref_1525_addr_0_ack_0 : boolean;
  signal ptr_deref_1525_load_0_req_0 : boolean;
  signal ptr_deref_1525_load_0_ack_0 : boolean;
  signal ptr_deref_1525_load_0_req_1 : boolean;
  signal ptr_deref_1525_load_0_ack_1 : boolean;
  signal ptr_deref_1525_gather_scatter_req_0 : boolean;
  signal ptr_deref_1525_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1529_base_resize_req_0 : boolean;
  signal ptr_deref_1529_base_resize_ack_0 : boolean;
  signal ptr_deref_1529_root_address_inst_req_0 : boolean;
  signal ptr_deref_1529_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1529_addr_0_req_0 : boolean;
  signal ptr_deref_1529_addr_0_ack_0 : boolean;
  signal ptr_deref_1529_load_0_req_0 : boolean;
  signal ptr_deref_1529_load_0_ack_0 : boolean;
  signal ptr_deref_1529_load_0_req_1 : boolean;
  signal ptr_deref_1529_load_0_ack_1 : boolean;
  signal ptr_deref_1529_gather_scatter_req_0 : boolean;
  signal ptr_deref_1529_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1533_base_resize_req_0 : boolean;
  signal ptr_deref_1533_base_resize_ack_0 : boolean;
  signal ptr_deref_1533_root_address_inst_req_0 : boolean;
  signal ptr_deref_1533_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1533_addr_0_req_0 : boolean;
  signal ptr_deref_1533_addr_0_ack_0 : boolean;
  signal ptr_deref_1533_load_0_req_0 : boolean;
  signal ptr_deref_1533_load_0_ack_0 : boolean;
  signal ptr_deref_1533_load_0_req_1 : boolean;
  signal ptr_deref_1533_load_0_ack_1 : boolean;
  signal ptr_deref_1533_gather_scatter_req_0 : boolean;
  signal ptr_deref_1533_gather_scatter_ack_0 : boolean;
  signal binary_1538_inst_req_0 : boolean;
  signal binary_1538_inst_ack_0 : boolean;
  signal binary_1538_inst_req_1 : boolean;
  signal binary_1538_inst_ack_1 : boolean;
  signal binary_1543_inst_req_0 : boolean;
  signal binary_1543_inst_ack_0 : boolean;
  signal binary_1543_inst_req_1 : boolean;
  signal binary_1543_inst_ack_1 : boolean;
  signal binary_1548_inst_req_0 : boolean;
  signal binary_1548_inst_ack_0 : boolean;
  signal binary_1548_inst_req_1 : boolean;
  signal binary_1548_inst_ack_1 : boolean;
  signal binary_1553_inst_req_0 : boolean;
  signal binary_1553_inst_ack_0 : boolean;
  signal binary_1553_inst_req_1 : boolean;
  signal binary_1553_inst_ack_1 : boolean;
  signal binary_1558_inst_req_0 : boolean;
  signal binary_1558_inst_ack_0 : boolean;
  signal binary_1558_inst_req_1 : boolean;
  signal binary_1558_inst_ack_1 : boolean;
  signal binary_1563_inst_req_0 : boolean;
  signal binary_1563_inst_ack_0 : boolean;
  signal binary_1563_inst_req_1 : boolean;
  signal binary_1563_inst_ack_1 : boolean;
  signal binary_1799_inst_req_1 : boolean;
  signal binary_1799_inst_ack_1 : boolean;
  signal binary_1819_inst_req_0 : boolean;
  signal binary_1568_inst_req_0 : boolean;
  signal binary_1568_inst_ack_0 : boolean;
  signal binary_1568_inst_req_1 : boolean;
  signal binary_1568_inst_ack_1 : boolean;
  signal ptr_deref_1976_root_address_inst_ack_0 : boolean;
  signal binary_1573_inst_req_0 : boolean;
  signal binary_1573_inst_ack_0 : boolean;
  signal binary_1573_inst_req_1 : boolean;
  signal binary_1573_inst_ack_1 : boolean;
  signal binary_1809_inst_req_0 : boolean;
  signal binary_1819_inst_ack_0 : boolean;
  signal binary_1809_inst_ack_0 : boolean;
  signal binary_1578_inst_req_0 : boolean;
  signal binary_1578_inst_ack_0 : boolean;
  signal binary_1578_inst_req_1 : boolean;
  signal binary_1578_inst_ack_1 : boolean;
  signal binary_1819_inst_ack_1 : boolean;
  signal binary_1809_inst_req_1 : boolean;
  signal binary_1809_inst_ack_1 : boolean;
  signal binary_1804_inst_req_0 : boolean;
  signal binary_1814_inst_req_0 : boolean;
  signal binary_1814_inst_ack_0 : boolean;
  signal binary_1804_inst_ack_0 : boolean;
  signal binary_1583_inst_req_0 : boolean;
  signal binary_1583_inst_ack_0 : boolean;
  signal binary_1583_inst_req_1 : boolean;
  signal binary_1583_inst_ack_1 : boolean;
  signal binary_1804_inst_req_1 : boolean;
  signal binary_1814_inst_req_1 : boolean;
  signal binary_1804_inst_ack_1 : boolean;
  signal binary_1814_inst_ack_1 : boolean;
  signal binary_1588_inst_req_0 : boolean;
  signal binary_1588_inst_ack_0 : boolean;
  signal binary_1588_inst_req_1 : boolean;
  signal binary_1588_inst_ack_1 : boolean;
  signal binary_1819_inst_req_1 : boolean;
  signal binary_1593_inst_req_0 : boolean;
  signal binary_1593_inst_ack_0 : boolean;
  signal binary_1593_inst_req_1 : boolean;
  signal binary_1593_inst_ack_1 : boolean;
  signal binary_1598_inst_req_0 : boolean;
  signal binary_1598_inst_ack_0 : boolean;
  signal binary_1598_inst_req_1 : boolean;
  signal binary_1598_inst_ack_1 : boolean;
  signal binary_1603_inst_req_0 : boolean;
  signal binary_1603_inst_ack_0 : boolean;
  signal binary_1603_inst_req_1 : boolean;
  signal binary_1603_inst_ack_1 : boolean;
  signal binary_1608_inst_req_0 : boolean;
  signal binary_1608_inst_ack_0 : boolean;
  signal binary_1608_inst_req_1 : boolean;
  signal binary_1608_inst_ack_1 : boolean;
  signal binary_1613_inst_req_0 : boolean;
  signal binary_1613_inst_ack_0 : boolean;
  signal binary_1613_inst_req_1 : boolean;
  signal binary_1613_inst_ack_1 : boolean;
  signal binary_1618_inst_req_0 : boolean;
  signal binary_1618_inst_ack_0 : boolean;
  signal binary_1618_inst_req_1 : boolean;
  signal binary_1618_inst_ack_1 : boolean;
  signal binary_1623_inst_req_0 : boolean;
  signal binary_1623_inst_ack_0 : boolean;
  signal binary_1623_inst_req_1 : boolean;
  signal binary_1623_inst_ack_1 : boolean;
  signal binary_1628_inst_req_0 : boolean;
  signal binary_1628_inst_ack_0 : boolean;
  signal binary_1628_inst_req_1 : boolean;
  signal binary_1628_inst_ack_1 : boolean;
  signal binary_1633_inst_req_0 : boolean;
  signal binary_1633_inst_ack_0 : boolean;
  signal binary_1668_inst_req_0 : boolean;
  signal binary_1668_inst_ack_0 : boolean;
  signal binary_1668_inst_req_1 : boolean;
  signal binary_1668_inst_ack_1 : boolean;
  signal binary_1673_inst_req_0 : boolean;
  signal binary_1673_inst_ack_0 : boolean;
  signal binary_1673_inst_req_1 : boolean;
  signal binary_1673_inst_ack_1 : boolean;
  signal binary_1678_inst_req_0 : boolean;
  signal binary_1678_inst_ack_0 : boolean;
  signal binary_1678_inst_req_1 : boolean;
  signal binary_1678_inst_ack_1 : boolean;
  signal binary_1683_inst_req_0 : boolean;
  signal binary_1683_inst_ack_0 : boolean;
  signal binary_1683_inst_req_1 : boolean;
  signal binary_1683_inst_ack_1 : boolean;
  signal binary_1688_inst_req_0 : boolean;
  signal binary_1688_inst_ack_0 : boolean;
  signal binary_1688_inst_req_1 : boolean;
  signal binary_1688_inst_ack_1 : boolean;
  signal binary_1693_inst_req_0 : boolean;
  signal binary_1693_inst_ack_0 : boolean;
  signal binary_1693_inst_req_1 : boolean;
  signal binary_1693_inst_ack_1 : boolean;
  signal ptr_deref_1980_root_address_inst_req_0 : boolean;
  signal ptr_deref_1697_base_resize_req_0 : boolean;
  signal ptr_deref_1697_base_resize_ack_0 : boolean;
  signal ptr_deref_1972_base_resize_req_0 : boolean;
  signal ptr_deref_1697_root_address_inst_req_0 : boolean;
  signal ptr_deref_1697_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1697_addr_0_req_0 : boolean;
  signal ptr_deref_1697_addr_0_ack_0 : boolean;
  signal ptr_deref_1972_base_resize_ack_0 : boolean;
  signal ptr_deref_1697_load_0_req_0 : boolean;
  signal ptr_deref_1697_load_0_ack_0 : boolean;
  signal ptr_deref_1697_load_0_req_1 : boolean;
  signal ptr_deref_1697_load_0_ack_1 : boolean;
  signal ptr_deref_1697_gather_scatter_req_0 : boolean;
  signal ptr_deref_1697_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1972_root_address_inst_req_0 : boolean;
  signal ptr_deref_1972_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1968_base_resize_req_0 : boolean;
  signal ptr_deref_1968_base_resize_ack_0 : boolean;
  signal ptr_deref_1701_base_resize_req_0 : boolean;
  signal ptr_deref_1701_base_resize_ack_0 : boolean;
  signal ptr_deref_1701_root_address_inst_req_0 : boolean;
  signal ptr_deref_1701_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1701_addr_0_req_0 : boolean;
  signal ptr_deref_1701_addr_0_ack_0 : boolean;
  signal ptr_deref_1972_addr_0_req_0 : boolean;
  signal ptr_deref_1701_load_0_req_0 : boolean;
  signal ptr_deref_1701_load_0_ack_0 : boolean;
  signal ptr_deref_1968_root_address_inst_req_0 : boolean;
  signal ptr_deref_1968_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1701_load_0_req_1 : boolean;
  signal ptr_deref_1701_load_0_ack_1 : boolean;
  signal ptr_deref_1701_gather_scatter_req_0 : boolean;
  signal ptr_deref_1701_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1980_store_0_req_1 : boolean;
  signal ptr_deref_1976_store_0_ack_1 : boolean;
  signal ptr_deref_1968_addr_0_req_0 : boolean;
  signal ptr_deref_1980_store_0_req_0 : boolean;
  signal ptr_deref_1968_addr_0_ack_0 : boolean;
  signal ptr_deref_1705_base_resize_req_0 : boolean;
  signal ptr_deref_1705_base_resize_ack_0 : boolean;
  signal ptr_deref_1705_root_address_inst_req_0 : boolean;
  signal ptr_deref_1705_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1980_gather_scatter_req_0 : boolean;
  signal ptr_deref_1972_addr_0_ack_0 : boolean;
  signal ptr_deref_1976_addr_0_req_0 : boolean;
  signal ptr_deref_1705_addr_0_req_0 : boolean;
  signal ptr_deref_1705_addr_0_ack_0 : boolean;
  signal ptr_deref_1968_gather_scatter_req_0 : boolean;
  signal ptr_deref_1705_load_0_req_0 : boolean;
  signal ptr_deref_1968_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1705_load_0_ack_0 : boolean;
  signal ptr_deref_1705_load_0_req_1 : boolean;
  signal ptr_deref_1705_load_0_ack_1 : boolean;
  signal ptr_deref_1705_gather_scatter_req_0 : boolean;
  signal ptr_deref_1705_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1976_store_0_ack_0 : boolean;
  signal ptr_deref_1980_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1968_store_0_req_0 : boolean;
  signal ptr_deref_1968_store_0_ack_0 : boolean;
  signal ptr_deref_1709_base_resize_req_0 : boolean;
  signal ptr_deref_1709_base_resize_ack_0 : boolean;
  signal ptr_deref_1980_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1709_root_address_inst_req_0 : boolean;
  signal ptr_deref_1709_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1972_gather_scatter_req_0 : boolean;
  signal ptr_deref_1709_addr_0_req_0 : boolean;
  signal ptr_deref_1709_addr_0_ack_0 : boolean;
  signal ptr_deref_1972_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1709_load_0_req_0 : boolean;
  signal ptr_deref_1709_load_0_ack_0 : boolean;
  signal ptr_deref_1709_load_0_req_1 : boolean;
  signal ptr_deref_1709_load_0_ack_1 : boolean;
  signal ptr_deref_1709_gather_scatter_req_0 : boolean;
  signal ptr_deref_1709_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1980_store_0_ack_0 : boolean;
  signal ptr_deref_1976_store_0_req_1 : boolean;
  signal ptr_deref_1976_store_0_req_0 : boolean;
  signal ptr_deref_1976_base_resize_ack_0 : boolean;
  signal ptr_deref_1976_addr_0_ack_0 : boolean;
  signal ptr_deref_1972_store_0_req_0 : boolean;
  signal ptr_deref_1968_store_0_req_1 : boolean;
  signal binary_1714_inst_req_0 : boolean;
  signal binary_1714_inst_ack_0 : boolean;
  signal binary_1714_inst_req_1 : boolean;
  signal binary_1714_inst_ack_1 : boolean;
  signal ptr_deref_1968_store_0_ack_1 : boolean;
  signal ptr_deref_1972_store_0_ack_0 : boolean;
  signal ptr_deref_1980_store_0_ack_1 : boolean;
  signal binary_1719_inst_req_0 : boolean;
  signal binary_1719_inst_ack_0 : boolean;
  signal binary_1719_inst_req_1 : boolean;
  signal binary_1719_inst_ack_1 : boolean;
  signal ptr_deref_1976_gather_scatter_req_0 : boolean;
  signal ptr_deref_1976_root_address_inst_req_0 : boolean;
  signal ptr_deref_1980_addr_0_req_0 : boolean;
  signal binary_1724_inst_req_0 : boolean;
  signal binary_1724_inst_ack_0 : boolean;
  signal binary_1724_inst_req_1 : boolean;
  signal binary_1724_inst_ack_1 : boolean;
  signal ptr_deref_1976_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1976_base_resize_req_0 : boolean;
  signal ptr_deref_1972_store_0_req_1 : boolean;
  signal binary_1729_inst_req_0 : boolean;
  signal binary_1729_inst_ack_0 : boolean;
  signal binary_1729_inst_req_1 : boolean;
  signal binary_1729_inst_ack_1 : boolean;
  signal binary_1734_inst_req_0 : boolean;
  signal binary_1734_inst_ack_0 : boolean;
  signal binary_1734_inst_req_1 : boolean;
  signal binary_1734_inst_ack_1 : boolean;
  signal binary_1739_inst_req_0 : boolean;
  signal binary_1739_inst_ack_0 : boolean;
  signal binary_1739_inst_req_1 : boolean;
  signal binary_1739_inst_ack_1 : boolean;
  signal binary_1744_inst_req_0 : boolean;
  signal binary_1744_inst_ack_0 : boolean;
  signal binary_1744_inst_req_1 : boolean;
  signal binary_1744_inst_ack_1 : boolean;
  signal binary_1749_inst_req_0 : boolean;
  signal binary_1749_inst_ack_0 : boolean;
  signal binary_1749_inst_req_1 : boolean;
  signal binary_1749_inst_ack_1 : boolean;
  signal binary_1754_inst_req_0 : boolean;
  signal binary_1754_inst_ack_0 : boolean;
  signal binary_1754_inst_req_1 : boolean;
  signal binary_1754_inst_ack_1 : boolean;
  signal binary_1759_inst_req_0 : boolean;
  signal binary_1759_inst_ack_0 : boolean;
  signal binary_1759_inst_req_1 : boolean;
  signal binary_1759_inst_ack_1 : boolean;
  signal binary_1764_inst_req_0 : boolean;
  signal binary_1764_inst_ack_0 : boolean;
  signal binary_1764_inst_req_1 : boolean;
  signal binary_1764_inst_ack_1 : boolean;
  signal binary_1769_inst_req_0 : boolean;
  signal binary_1769_inst_ack_0 : boolean;
  signal binary_1769_inst_req_1 : boolean;
  signal binary_1769_inst_ack_1 : boolean;
  signal binary_1774_inst_req_0 : boolean;
  signal binary_1774_inst_ack_0 : boolean;
  signal binary_1774_inst_req_1 : boolean;
  signal binary_1774_inst_ack_1 : boolean;
  signal binary_1779_inst_req_0 : boolean;
  signal binary_1779_inst_ack_0 : boolean;
  signal binary_1779_inst_req_1 : boolean;
  signal binary_1779_inst_ack_1 : boolean;
  signal binary_1784_inst_req_0 : boolean;
  signal binary_1784_inst_ack_0 : boolean;
  signal binary_1784_inst_req_1 : boolean;
  signal binary_1784_inst_ack_1 : boolean;
  signal ptr_deref_1980_base_resize_ack_0 : boolean;
  signal binary_1789_inst_req_0 : boolean;
  signal binary_1789_inst_ack_0 : boolean;
  signal binary_1789_inst_req_1 : boolean;
  signal binary_1789_inst_ack_1 : boolean;
  signal ptr_deref_1980_base_resize_req_0 : boolean;
  signal binary_1794_inst_req_0 : boolean;
  signal binary_1794_inst_ack_0 : boolean;
  signal binary_1794_inst_req_1 : boolean;
  signal binary_1794_inst_ack_1 : boolean;
  signal binary_1799_inst_req_0 : boolean;
  signal binary_1799_inst_ack_0 : boolean;
  signal binary_1824_inst_req_0 : boolean;
  signal binary_1824_inst_ack_0 : boolean;
  signal binary_1824_inst_req_1 : boolean;
  signal binary_1824_inst_ack_1 : boolean;
  signal binary_1829_inst_req_0 : boolean;
  signal binary_1829_inst_ack_0 : boolean;
  signal binary_1829_inst_req_1 : boolean;
  signal binary_1829_inst_ack_1 : boolean;
  signal binary_1834_inst_req_0 : boolean;
  signal binary_1834_inst_ack_0 : boolean;
  signal binary_1834_inst_req_1 : boolean;
  signal binary_1834_inst_ack_1 : boolean;
  signal ptr_deref_1972_store_0_ack_1 : boolean;
  signal phi_stmt_813_req_1 : boolean;
  signal binary_1839_inst_req_0 : boolean;
  signal binary_1839_inst_ack_0 : boolean;
  signal binary_1839_inst_req_1 : boolean;
  signal binary_1839_inst_ack_1 : boolean;
  signal type_cast_847_inst_req_0 : boolean;
  signal type_cast_847_inst_ack_0 : boolean;
  signal binary_1844_inst_req_0 : boolean;
  signal binary_1844_inst_ack_0 : boolean;
  signal type_cast_777_inst_req_0 : boolean;
  signal binary_1844_inst_req_1 : boolean;
  signal binary_1844_inst_ack_1 : boolean;
  signal type_cast_777_inst_ack_0 : boolean;
  signal binary_1849_inst_req_0 : boolean;
  signal phi_stmt_771_req_1 : boolean;
  signal binary_1849_inst_ack_0 : boolean;
  signal binary_1849_inst_req_1 : boolean;
  signal binary_1849_inst_ack_1 : boolean;
  signal type_cast_826_inst_req_0 : boolean;
  signal type_cast_826_inst_ack_0 : boolean;
  signal phi_stmt_820_req_1 : boolean;
  signal phi_stmt_841_req_1 : boolean;
  signal binary_1854_inst_req_0 : boolean;
  signal binary_1854_inst_ack_0 : boolean;
  signal binary_1854_inst_req_1 : boolean;
  signal binary_1854_inst_ack_1 : boolean;
  signal type_cast_784_inst_req_0 : boolean;
  signal type_cast_784_inst_ack_0 : boolean;
  signal phi_stmt_778_req_0 : boolean;
  signal phi_stmt_778_req_1 : boolean;
  signal binary_1859_inst_req_0 : boolean;
  signal binary_1859_inst_ack_0 : boolean;
  signal binary_1859_inst_req_1 : boolean;
  signal binary_1859_inst_ack_1 : boolean;
  signal type_cast_833_inst_req_0 : boolean;
  signal type_cast_833_inst_ack_0 : boolean;
  signal phi_stmt_827_req_1 : boolean;
  signal binary_1864_inst_req_0 : boolean;
  signal binary_1864_inst_ack_0 : boolean;
  signal binary_1864_inst_req_1 : boolean;
  signal binary_1864_inst_ack_1 : boolean;
  signal type_cast_791_inst_req_0 : boolean;
  signal type_cast_791_inst_ack_0 : boolean;
  signal phi_stmt_785_req_1 : boolean;
  signal phi_stmt_771_req_0 : boolean;
  signal binary_1869_inst_req_0 : boolean;
  signal binary_1869_inst_ack_0 : boolean;
  signal binary_1869_inst_req_1 : boolean;
  signal binary_1869_inst_ack_1 : boolean;
  signal type_cast_840_inst_req_0 : boolean;
  signal type_cast_840_inst_ack_0 : boolean;
  signal type_cast_798_inst_req_0 : boolean;
  signal type_cast_798_inst_ack_0 : boolean;
  signal type_cast_861_inst_req_0 : boolean;
  signal phi_stmt_792_req_1 : boolean;
  signal binary_1875_inst_req_0 : boolean;
  signal binary_1875_inst_ack_0 : boolean;
  signal binary_1875_inst_req_1 : boolean;
  signal binary_1875_inst_ack_1 : boolean;
  signal phi_stmt_834_req_1 : boolean;
  signal type_cast_861_inst_ack_0 : boolean;
  signal phi_stmt_855_req_1 : boolean;
  signal phi_stmt_750_req_0 : boolean;
  signal binary_1881_inst_req_0 : boolean;
  signal binary_1881_inst_ack_0 : boolean;
  signal binary_1881_inst_req_1 : boolean;
  signal binary_1881_inst_ack_1 : boolean;
  signal if_stmt_1883_branch_req_0 : boolean;
  signal if_stmt_1883_branch_ack_1 : boolean;
  signal if_stmt_1883_branch_ack_0 : boolean;
  signal ptr_deref_1956_base_resize_req_0 : boolean;
  signal ptr_deref_1956_base_resize_ack_0 : boolean;
  signal ptr_deref_1956_root_address_inst_req_0 : boolean;
  signal ptr_deref_1956_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1956_addr_0_req_0 : boolean;
  signal ptr_deref_1956_addr_0_ack_0 : boolean;
  signal ptr_deref_1956_gather_scatter_req_0 : boolean;
  signal ptr_deref_1956_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1956_store_0_req_0 : boolean;
  signal ptr_deref_1956_store_0_ack_0 : boolean;
  signal ptr_deref_1956_store_0_req_1 : boolean;
  signal ptr_deref_1956_store_0_ack_1 : boolean;
  signal ptr_deref_1980_addr_0_ack_0 : boolean;
  signal ptr_deref_1960_base_resize_req_0 : boolean;
  signal ptr_deref_1960_base_resize_ack_0 : boolean;
  signal ptr_deref_1960_root_address_inst_req_0 : boolean;
  signal ptr_deref_1960_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1960_addr_0_req_0 : boolean;
  signal ptr_deref_1960_addr_0_ack_0 : boolean;
  signal ptr_deref_1960_gather_scatter_req_0 : boolean;
  signal ptr_deref_1960_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1960_store_0_req_0 : boolean;
  signal ptr_deref_1960_store_0_ack_0 : boolean;
  signal ptr_deref_1960_store_0_req_1 : boolean;
  signal ptr_deref_1960_store_0_ack_1 : boolean;
  signal ptr_deref_1964_base_resize_req_0 : boolean;
  signal ptr_deref_1964_base_resize_ack_0 : boolean;
  signal ptr_deref_1964_root_address_inst_req_0 : boolean;
  signal ptr_deref_1964_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1964_addr_0_req_0 : boolean;
  signal ptr_deref_1964_addr_0_ack_0 : boolean;
  signal ptr_deref_1964_gather_scatter_req_0 : boolean;
  signal ptr_deref_1964_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1964_store_0_req_0 : boolean;
  signal ptr_deref_1964_store_0_ack_0 : boolean;
  signal ptr_deref_1964_store_0_req_1 : boolean;
  signal ptr_deref_1964_store_0_ack_1 : boolean;
  signal ptr_deref_1984_base_resize_req_0 : boolean;
  signal ptr_deref_1984_base_resize_ack_0 : boolean;
  signal ptr_deref_1984_root_address_inst_req_0 : boolean;
  signal ptr_deref_1984_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1984_addr_0_req_0 : boolean;
  signal ptr_deref_1984_addr_0_ack_0 : boolean;
  signal ptr_deref_1984_gather_scatter_req_0 : boolean;
  signal ptr_deref_1984_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1984_store_0_req_0 : boolean;
  signal ptr_deref_1984_store_0_ack_0 : boolean;
  signal ptr_deref_1984_store_0_req_1 : boolean;
  signal ptr_deref_1984_store_0_ack_1 : boolean;
  signal ptr_deref_1988_base_resize_req_0 : boolean;
  signal ptr_deref_1988_base_resize_ack_0 : boolean;
  signal ptr_deref_1988_root_address_inst_req_0 : boolean;
  signal ptr_deref_1988_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1988_addr_0_req_0 : boolean;
  signal ptr_deref_1988_addr_0_ack_0 : boolean;
  signal ptr_deref_1988_gather_scatter_req_0 : boolean;
  signal ptr_deref_1988_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1988_store_0_req_0 : boolean;
  signal ptr_deref_1988_store_0_ack_0 : boolean;
  signal ptr_deref_1988_store_0_req_1 : boolean;
  signal ptr_deref_1988_store_0_ack_1 : boolean;
  signal ptr_deref_1992_base_resize_req_0 : boolean;
  signal ptr_deref_1992_base_resize_ack_0 : boolean;
  signal ptr_deref_1992_root_address_inst_req_0 : boolean;
  signal ptr_deref_1992_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1992_addr_0_req_0 : boolean;
  signal ptr_deref_1992_addr_0_ack_0 : boolean;
  signal ptr_deref_1992_gather_scatter_req_0 : boolean;
  signal ptr_deref_1992_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1992_store_0_req_0 : boolean;
  signal ptr_deref_1992_store_0_ack_0 : boolean;
  signal ptr_deref_1992_store_0_req_1 : boolean;
  signal ptr_deref_1992_store_0_ack_1 : boolean;
  signal ptr_deref_1996_base_resize_req_0 : boolean;
  signal ptr_deref_1996_base_resize_ack_0 : boolean;
  signal ptr_deref_1996_root_address_inst_req_0 : boolean;
  signal ptr_deref_1996_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1996_addr_0_req_0 : boolean;
  signal ptr_deref_1996_addr_0_ack_0 : boolean;
  signal ptr_deref_1996_gather_scatter_req_0 : boolean;
  signal ptr_deref_1996_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1996_store_0_req_0 : boolean;
  signal ptr_deref_1996_store_0_ack_0 : boolean;
  signal ptr_deref_1996_store_0_req_1 : boolean;
  signal ptr_deref_1996_store_0_ack_1 : boolean;
  signal ptr_deref_2000_base_resize_req_0 : boolean;
  signal ptr_deref_2000_base_resize_ack_0 : boolean;
  signal ptr_deref_2000_root_address_inst_req_0 : boolean;
  signal ptr_deref_2000_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2000_addr_0_req_0 : boolean;
  signal ptr_deref_2000_addr_0_ack_0 : boolean;
  signal ptr_deref_2000_gather_scatter_req_0 : boolean;
  signal ptr_deref_2000_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2000_store_0_req_0 : boolean;
  signal ptr_deref_2000_store_0_ack_0 : boolean;
  signal ptr_deref_2000_store_0_req_1 : boolean;
  signal ptr_deref_2000_store_0_ack_1 : boolean;
  signal type_cast_819_inst_ack_0 : boolean;
  signal phi_stmt_848_req_1 : boolean;
  signal type_cast_819_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal phi_stmt_743_req_0 : boolean;
  signal phi_stmt_792_req_0 : boolean;
  signal phi_stmt_764_req_1 : boolean;
  signal type_cast_770_inst_ack_0 : boolean;
  signal type_cast_770_inst_req_0 : boolean;
  signal phi_stmt_799_req_0 : boolean;
  signal phi_stmt_757_req_1 : boolean;
  signal type_cast_763_inst_ack_0 : boolean;
  signal type_cast_763_inst_req_0 : boolean;
  signal ptr_deref_2004_base_resize_req_0 : boolean;
  signal ptr_deref_2004_base_resize_ack_0 : boolean;
  signal ptr_deref_2004_root_address_inst_req_0 : boolean;
  signal ptr_deref_2004_root_address_inst_ack_0 : boolean;
  signal phi_stmt_806_req_0 : boolean;
  signal ptr_deref_2004_addr_0_req_0 : boolean;
  signal phi_stmt_750_req_1 : boolean;
  signal ptr_deref_2004_addr_0_ack_0 : boolean;
  signal type_cast_756_inst_ack_0 : boolean;
  signal ptr_deref_2004_gather_scatter_req_0 : boolean;
  signal type_cast_756_inst_req_0 : boolean;
  signal ptr_deref_2004_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2004_store_0_req_0 : boolean;
  signal ptr_deref_2004_store_0_ack_0 : boolean;
  signal phi_stmt_757_req_0 : boolean;
  signal ptr_deref_2004_store_0_req_1 : boolean;
  signal ptr_deref_2004_store_0_ack_1 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal phi_stmt_806_req_1 : boolean;
  signal type_cast_812_inst_ack_0 : boolean;
  signal phi_stmt_743_req_1 : boolean;
  signal type_cast_749_inst_ack_0 : boolean;
  signal phi_stmt_785_req_0 : boolean;
  signal type_cast_812_inst_req_0 : boolean;
  signal type_cast_749_inst_req_0 : boolean;
  signal ptr_deref_2008_base_resize_req_0 : boolean;
  signal phi_stmt_589_ack_0 : boolean;
  signal ptr_deref_2008_base_resize_ack_0 : boolean;
  signal phi_stmt_799_req_1 : boolean;
  signal ptr_deref_2008_root_address_inst_req_0 : boolean;
  signal ptr_deref_2008_root_address_inst_ack_0 : boolean;
  signal type_cast_805_inst_ack_0 : boolean;
  signal type_cast_805_inst_req_0 : boolean;
  signal ptr_deref_2008_addr_0_req_0 : boolean;
  signal ptr_deref_2008_addr_0_ack_0 : boolean;
  signal ptr_deref_2008_gather_scatter_req_0 : boolean;
  signal ptr_deref_2008_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2008_store_0_req_0 : boolean;
  signal ptr_deref_2008_store_0_ack_0 : boolean;
  signal ptr_deref_2008_store_0_req_1 : boolean;
  signal ptr_deref_2008_store_0_ack_1 : boolean;
  signal ptr_deref_2012_base_resize_req_0 : boolean;
  signal ptr_deref_2012_base_resize_ack_0 : boolean;
  signal ptr_deref_2012_root_address_inst_req_0 : boolean;
  signal ptr_deref_2012_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2012_addr_0_req_0 : boolean;
  signal ptr_deref_2012_addr_0_ack_0 : boolean;
  signal ptr_deref_2012_gather_scatter_req_0 : boolean;
  signal ptr_deref_2012_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2012_store_0_req_0 : boolean;
  signal ptr_deref_2012_store_0_ack_0 : boolean;
  signal ptr_deref_2012_store_0_req_1 : boolean;
  signal ptr_deref_2012_store_0_ack_1 : boolean;
  signal ptr_deref_2016_base_resize_req_0 : boolean;
  signal ptr_deref_2016_base_resize_ack_0 : boolean;
  signal ptr_deref_2016_root_address_inst_req_0 : boolean;
  signal ptr_deref_2016_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2016_addr_0_req_0 : boolean;
  signal ptr_deref_2016_addr_0_ack_0 : boolean;
  signal ptr_deref_2016_gather_scatter_req_0 : boolean;
  signal ptr_deref_2016_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2016_store_0_req_0 : boolean;
  signal ptr_deref_2016_store_0_ack_0 : boolean;
  signal ptr_deref_2016_store_0_req_1 : boolean;
  signal ptr_deref_2016_store_0_ack_1 : boolean;
  signal binary_2023_inst_req_0 : boolean;
  signal binary_2023_inst_ack_0 : boolean;
  signal binary_2023_inst_req_1 : boolean;
  signal binary_2023_inst_ack_1 : boolean;
  signal binary_2029_inst_req_0 : boolean;
  signal binary_2029_inst_ack_0 : boolean;
  signal binary_2029_inst_req_1 : boolean;
  signal binary_2029_inst_ack_1 : boolean;
  signal if_stmt_2031_branch_req_0 : boolean;
  signal if_stmt_2031_branch_ack_1 : boolean;
  signal if_stmt_2031_branch_ack_0 : boolean;
  signal binary_2042_inst_req_0 : boolean;
  signal binary_2042_inst_ack_0 : boolean;
  signal binary_2042_inst_req_1 : boolean;
  signal binary_2042_inst_ack_1 : boolean;
  signal binary_2048_inst_req_0 : boolean;
  signal binary_2048_inst_ack_0 : boolean;
  signal binary_2048_inst_req_1 : boolean;
  signal binary_2048_inst_ack_1 : boolean;
  signal if_stmt_2050_branch_req_0 : boolean;
  signal if_stmt_2050_branch_ack_1 : boolean;
  signal if_stmt_2050_branch_ack_0 : boolean;
  signal phi_stmt_555_req_0 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal phi_stmt_555_req_1 : boolean;
  signal phi_stmt_555_ack_0 : boolean;
  signal phi_stmt_589_req_0 : boolean;
  signal type_cast_595_inst_req_0 : boolean;
  signal type_cast_595_inst_ack_0 : boolean;
  signal phi_stmt_589_req_1 : boolean;
  signal phi_stmt_813_req_0 : boolean;
  signal phi_stmt_820_req_0 : boolean;
  signal phi_stmt_827_req_0 : boolean;
  signal phi_stmt_834_req_0 : boolean;
  signal phi_stmt_841_req_0 : boolean;
  signal phi_stmt_848_req_0 : boolean;
  signal phi_stmt_855_req_0 : boolean;
  signal phi_stmt_743_ack_0 : boolean;
  signal phi_stmt_750_ack_0 : boolean;
  signal phi_stmt_757_ack_0 : boolean;
  signal phi_stmt_764_ack_0 : boolean;
  signal phi_stmt_771_ack_0 : boolean;
  signal phi_stmt_778_ack_0 : boolean;
  signal phi_stmt_785_ack_0 : boolean;
  signal phi_stmt_792_ack_0 : boolean;
  signal phi_stmt_799_ack_0 : boolean;
  signal phi_stmt_806_ack_0 : boolean;
  signal phi_stmt_813_ack_0 : boolean;
  signal phi_stmt_820_ack_0 : boolean;
  signal phi_stmt_827_ack_0 : boolean;
  signal phi_stmt_834_ack_0 : boolean;
  signal phi_stmt_841_ack_0 : boolean;
  signal phi_stmt_848_ack_0 : boolean;
  signal phi_stmt_855_ack_0 : boolean;
  signal type_cast_1893_inst_req_0 : boolean;
  signal type_cast_1893_inst_ack_0 : boolean;
  signal phi_stmt_1890_req_0 : boolean;
  signal type_cast_1897_inst_req_0 : boolean;
  signal type_cast_1897_inst_ack_0 : boolean;
  signal phi_stmt_1894_req_0 : boolean;
  signal type_cast_1901_inst_req_0 : boolean;
  signal type_cast_1901_inst_ack_0 : boolean;
  signal phi_stmt_1898_req_0 : boolean;
  signal type_cast_1905_inst_req_0 : boolean;
  signal type_cast_1905_inst_ack_0 : boolean;
  signal phi_stmt_1902_req_0 : boolean;
  signal type_cast_1909_inst_req_0 : boolean;
  signal type_cast_1909_inst_ack_0 : boolean;
  signal phi_stmt_1906_req_0 : boolean;
  signal type_cast_1913_inst_req_0 : boolean;
  signal type_cast_1913_inst_ack_0 : boolean;
  signal phi_stmt_1910_req_0 : boolean;
  signal type_cast_1917_inst_req_0 : boolean;
  signal type_cast_1917_inst_ack_0 : boolean;
  signal phi_stmt_1914_req_0 : boolean;
  signal type_cast_1921_inst_req_0 : boolean;
  signal type_cast_1921_inst_ack_0 : boolean;
  signal phi_stmt_1918_req_0 : boolean;
  signal type_cast_1925_inst_req_0 : boolean;
  signal type_cast_1925_inst_ack_0 : boolean;
  signal phi_stmt_1922_req_0 : boolean;
  signal type_cast_1929_inst_req_0 : boolean;
  signal type_cast_1929_inst_ack_0 : boolean;
  signal phi_stmt_1926_req_0 : boolean;
  signal type_cast_1933_inst_req_0 : boolean;
  signal type_cast_1933_inst_ack_0 : boolean;
  signal phi_stmt_1930_req_0 : boolean;
  signal type_cast_1937_inst_req_0 : boolean;
  signal type_cast_1937_inst_ack_0 : boolean;
  signal phi_stmt_1934_req_0 : boolean;
  signal type_cast_1941_inst_req_0 : boolean;
  signal type_cast_1941_inst_ack_0 : boolean;
  signal phi_stmt_1938_req_0 : boolean;
  signal type_cast_1945_inst_req_0 : boolean;
  signal type_cast_1945_inst_ack_0 : boolean;
  signal phi_stmt_1942_req_0 : boolean;
  signal type_cast_1949_inst_req_0 : boolean;
  signal type_cast_1949_inst_ack_0 : boolean;
  signal phi_stmt_1946_req_0 : boolean;
  signal type_cast_1953_inst_req_0 : boolean;
  signal type_cast_1953_inst_ack_0 : boolean;
  signal phi_stmt_1950_req_0 : boolean;
  signal phi_stmt_1890_ack_0 : boolean;
  signal phi_stmt_1894_ack_0 : boolean;
  signal phi_stmt_1898_ack_0 : boolean;
  signal phi_stmt_1902_ack_0 : boolean;
  signal phi_stmt_1906_ack_0 : boolean;
  signal phi_stmt_1910_ack_0 : boolean;
  signal phi_stmt_1914_ack_0 : boolean;
  signal phi_stmt_1918_ack_0 : boolean;
  signal phi_stmt_1922_ack_0 : boolean;
  signal phi_stmt_1926_ack_0 : boolean;
  signal phi_stmt_1930_ack_0 : boolean;
  signal phi_stmt_1934_ack_0 : boolean;
  signal phi_stmt_1938_ack_0 : boolean;
  signal phi_stmt_1942_ack_0 : boolean;
  signal phi_stmt_1946_ack_0 : boolean;
  signal phi_stmt_1950_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  mmultiply_base_CP_1311: Block -- control-path 
    signal cp_elements: BooleanArray(2777 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(8);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(8), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  output  bypass 
    -- predecessors 
    -- successors 2637 
    -- members (15) 
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36
      -- 	branch_block_stmt_552/branch_block_stmt_552__entry__
      -- 	branch_block_stmt_552/$entry
      -- 	$entry
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/$entry
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/$exit
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/$entry
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/$exit
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/$entry
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/$exit
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/req
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/ack
      -- 	branch_block_stmt_552/bbx_xnph39_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_req
      -- 
    phi_stmt_555_req_10169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => phi_stmt_555_req_0); -- 
    -- CP-element group 1 transition  place  output  bypass 
    -- predecessors 36 
    -- successors 2641 
    -- members (13) 
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586__exit__
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/$entry
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/$exit
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/$entry
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/$exit
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/$entry
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/$exit
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/req
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/ack
      -- 	branch_block_stmt_552/bbx_xnph36_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_req
      -- 
    cp_elements(1) <= cp_elements(36);
    phi_stmt_589_req_10204_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => phi_stmt_589_req_0); -- 
    -- CP-element group 2 place  bypass 
    -- predecessors 366 
    -- successors 2680 
    -- members (2) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740__exit__
      -- 
    cp_elements(2) <= cp_elements(366);
    -- CP-element group 3 place  bypass 
    -- predecessors 2718 
    -- successors 367 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882__entry__
      -- 	branch_block_stmt_552/merge_stmt_742__exit__
      -- 
    cp_elements(3) <= cp_elements(2718);
    -- CP-element group 4 branch  place  bypass 
    -- predecessors 2341 
    -- successors 2342 2345 
    -- members (2) 
      -- 	branch_block_stmt_552/if_stmt_1883__entry__
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882__exit__
      -- 
    cp_elements(4) <= cp_elements(2341);
    -- CP-element group 5 merge  place  bypass 
    -- predecessors 2720 2773 
    -- successors 2351 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030__entry__
      -- 	branch_block_stmt_552/merge_stmt_1889__exit__
      -- 
    cp_elements(5) <= OrReduce(cp_elements(2720) & cp_elements(2773));
    -- CP-element group 6 branch  place  bypass 
    -- predecessors 2605 
    -- successors 2606 2609 
    -- members (2) 
      -- 	branch_block_stmt_552/if_stmt_2031__entry__
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030__exit__
      -- 
    cp_elements(6) <= cp_elements(2605);
    -- CP-element group 7 merge  fork  transition  place  no-bypass 
    -- predecessors 2612 2775 
    -- successors 2615 2617 
    -- members (7) 
      -- 	branch_block_stmt_552/merge_stmt_2037__exit__
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049__entry__
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/$entry
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_trigger_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/simple_obj_ref_2039_trigger_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/simple_obj_ref_2039_active_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/simple_obj_ref_2039_completed_
      -- 
    cp_elements(7) <= OrReduce(cp_elements(2612) & cp_elements(2775));
    -- CP-element group 8 merge  transition  place  bypass 
    -- predecessors 2633 2777 
    -- successors 
    -- members (12) 
      -- 	branch_block_stmt_552/merge_stmt_2058__exit__
      -- 	branch_block_stmt_552/merge_stmt_2056__exit__
      -- 	branch_block_stmt_552/return__
      -- 	branch_block_stmt_552/branch_block_stmt_552__exit__
      -- 	branch_block_stmt_552/$exit
      -- 	$exit
      -- 	branch_block_stmt_552/merge_stmt_2058_PhiReqMerge
      -- 	branch_block_stmt_552/return___PhiReq/$entry
      -- 	branch_block_stmt_552/return___PhiReq/$exit
      -- 	branch_block_stmt_552/merge_stmt_2058_PhiAck/$entry
      -- 	branch_block_stmt_552/merge_stmt_2058_PhiAck/$exit
      -- 	branch_block_stmt_552/merge_stmt_2058_PhiAck/dummy
      -- 
    cp_elements(8) <= OrReduce(cp_elements(2633) & cp_elements(2777));
    -- CP-element group 9 join  fork  transition  bypass 
    -- predecessors 12 2639 
    -- successors 10 13 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_active_
      -- 
    cpelement_group_9 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(12);
      predecessors(1) <= cp_elements(2639);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(9)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(9),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 10 join  fork  transition  bypass 
    -- predecessors 9 14 
    -- successors 17 24 31 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_568_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_568_active_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_568_trigger_
      -- 
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(9);
      predecessors(1) <= cp_elements(14);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(10)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 11 transition  output  bypass 
    -- predecessors 2639 
    -- successors 12 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Sample/$entry
      -- 
    cp_elements(11) <= cp_elements(2639);
    rr_1364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => binary_567_inst_req_0); -- 
    -- CP-element group 12 transition  input  no-bypass 
    -- predecessors 11 
    -- successors 9 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Sample/$exit
      -- 
    ra_1365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_567_inst_ack_0, ack => cp_elements(12)); -- 
    -- CP-element group 13 transition  output  bypass 
    -- predecessors 9 
    -- successors 14 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Update/$entry
      -- 
    cp_elements(13) <= cp_elements(9);
    cr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => binary_567_inst_req_1); -- 
    -- CP-element group 14 transition  input  no-bypass 
    -- predecessors 13 
    -- successors 10 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_complete_Update/$exit
      -- 
    ca_1370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_567_inst_ack_1, ack => cp_elements(14)); -- 
    -- CP-element group 15 join  fork  transition  no-bypass 
    -- predecessors 17 19 
    -- successors 16 20 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_active_
      -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(17);
      predecessors(1) <= cp_elements(19);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(15)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 16 join  transition  no-bypass 
    -- predecessors 15 21 
    -- successors 36 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_574_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_574_active_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_574_trigger_
      -- 
    cpelement_group_16 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(15);
      predecessors(1) <= cp_elements(21);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(16)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(16),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 17 fork  transition  bypass 
    -- predecessors 10 
    -- successors 15 18 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_570_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_570_active_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_570_trigger_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_trigger_
      -- 
    cp_elements(17) <= cp_elements(10);
    -- CP-element group 18 transition  output  bypass 
    -- predecessors 17 
    -- successors 19 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Sample/$entry
      -- 
    cp_elements(18) <= cp_elements(17);
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_573_inst_req_0); -- 
    -- CP-element group 19 transition  input  no-bypass 
    -- predecessors 18 
    -- successors 15 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Sample/$exit
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_573_inst_ack_0, ack => cp_elements(19)); -- 
    -- CP-element group 20 transition  output  bypass 
    -- predecessors 15 
    -- successors 21 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Update/$entry
      -- 
    cp_elements(20) <= cp_elements(15);
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => binary_573_inst_req_1); -- 
    -- CP-element group 21 transition  input  no-bypass 
    -- predecessors 20 
    -- successors 16 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_573_complete_Update/$exit
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_573_inst_ack_1, ack => cp_elements(21)); -- 
    -- CP-element group 22 join  fork  transition  no-bypass 
    -- predecessors 24 26 
    -- successors 23 27 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_active_
      -- 
    cpelement_group_22 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(24);
      predecessors(1) <= cp_elements(26);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(22)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(22),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 23 join  transition  no-bypass 
    -- predecessors 22 28 
    -- successors 36 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_580_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_580_active_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_580_trigger_
      -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(22);
      predecessors(1) <= cp_elements(28);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(23)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 24 fork  transition  bypass 
    -- predecessors 10 
    -- successors 22 25 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_576_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_576_active_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_576_trigger_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_trigger_
      -- 
    cp_elements(24) <= cp_elements(10);
    -- CP-element group 25 transition  output  bypass 
    -- predecessors 24 
    -- successors 26 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Sample/$entry
      -- 
    cp_elements(25) <= cp_elements(24);
    rr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => binary_579_inst_req_0); -- 
    -- CP-element group 26 transition  input  no-bypass 
    -- predecessors 25 
    -- successors 22 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Sample/$exit
      -- 
    ra_1403_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_579_inst_ack_0, ack => cp_elements(26)); -- 
    -- CP-element group 27 transition  output  bypass 
    -- predecessors 22 
    -- successors 28 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Update/$entry
      -- 
    cp_elements(27) <= cp_elements(22);
    cr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => binary_579_inst_req_1); -- 
    -- CP-element group 28 transition  input  no-bypass 
    -- predecessors 27 
    -- successors 23 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_579_complete_Update/ca
      -- 
    ca_1408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_579_inst_ack_1, ack => cp_elements(28)); -- 
    -- CP-element group 29 join  fork  transition  no-bypass 
    -- predecessors 31 33 
    -- successors 30 34 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_active_
      -- 
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(31);
      predecessors(1) <= cp_elements(33);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(29)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 30 join  transition  no-bypass 
    -- predecessors 29 35 
    -- successors 36 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_586_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_586_active_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/assign_stmt_586_trigger_
      -- 
    cpelement_group_30 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(29);
      predecessors(1) <= cp_elements(35);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(30)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(30),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 31 fork  transition  bypass 
    -- predecessors 10 
    -- successors 29 32 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_582_trigger_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_trigger_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_582_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_582_active_
      -- 
    cp_elements(31) <= cp_elements(10);
    -- CP-element group 32 transition  output  bypass 
    -- predecessors 31 
    -- successors 33 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Sample/$entry
      -- 
    cp_elements(32) <= cp_elements(31);
    rr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => binary_585_inst_req_0); -- 
    -- CP-element group 33 transition  input  no-bypass 
    -- predecessors 32 
    -- successors 29 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Sample/$exit
      -- 
    ra_1422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_585_inst_ack_0, ack => cp_elements(33)); -- 
    -- CP-element group 34 transition  output  bypass 
    -- predecessors 29 
    -- successors 35 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Update/cr
      -- 
    cp_elements(34) <= cp_elements(29);
    cr_1426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => binary_585_inst_req_1); -- 
    -- CP-element group 35 transition  input  no-bypass 
    -- predecessors 34 
    -- successors 30 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_585_complete_Update/ca
      -- 
    ca_1427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_585_inst_ack_1, ack => cp_elements(35)); -- 
    -- CP-element group 36 join  transition  bypass 
    -- predecessors 16 23 30 
    -- successors 1 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/$exit
      -- 
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(16);
      predecessors(1) <= cp_elements(23);
      predecessors(2) <= cp_elements(30);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(36)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 37 fork  transition  bypass 
    -- predecessors 2643 
    -- successors 40 45 49 69 73 93 97 110 114 127 131 144 148 168 172 185 189 202 206 219 223 236 240 253 257 270 274 287 291 304 308 321 325 340 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/$entry
      -- 
    cp_elements(37) <= cp_elements(2643);
    -- CP-element group 38 join  fork  transition  bypass 
    -- predecessors 40 42 
    -- successors 39 43 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_active_
      -- 
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(40);
      predecessors(1) <= cp_elements(42);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(38)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 39 join  fork  transition  no-bypass 
    -- predecessors 38 44 
    -- successors 53 64 88 118 163 193 261 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_602_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_602_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_602_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_completed_
      -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(38);
      predecessors(1) <= cp_elements(44);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(39)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 40 fork  transition  bypass 
    -- predecessors 37 
    -- successors 38 41 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_598_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_598_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_598_trigger_
      -- 
    cp_elements(40) <= cp_elements(37);
    -- CP-element group 41 transition  output  bypass 
    -- predecessors 40 
    -- successors 42 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Sample/rr
      -- 
    cp_elements(41) <= cp_elements(40);
    rr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => binary_601_inst_req_0); -- 
    -- CP-element group 42 transition  input  no-bypass 
    -- predecessors 41 
    -- successors 38 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Sample/$exit
      -- 
    ra_1444_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_601_inst_ack_0, ack => cp_elements(42)); -- 
    -- CP-element group 43 transition  output  bypass 
    -- predecessors 38 
    -- successors 44 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Update/$entry
      -- 
    cp_elements(43) <= cp_elements(38);
    cr_1448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => binary_601_inst_req_1); -- 
    -- CP-element group 44 transition  input  no-bypass 
    -- predecessors 43 
    -- successors 39 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_601_complete_Update/ca
      -- 
    ca_1449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_601_inst_ack_1, ack => cp_elements(44)); -- 
    -- CP-element group 45 transition  bypass 
    -- predecessors 37 
    -- successors 46 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_607_trigger_
      -- 
    cp_elements(45) <= cp_elements(37);
    -- CP-element group 46 join  fork  transition  bypass 
    -- predecessors 45 59 
    -- successors 47 60 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_607_active_
      -- 
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(45);
      predecessors(1) <= cp_elements(59);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(46)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 47 join  transition  no-bypass 
    -- predecessors 46 61 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_608_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_608_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_607_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_608_completed_
      -- 
    cpelement_group_47 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(46);
      predecessors(1) <= cp_elements(61);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(47)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(47),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 48 join  transition  output  bypass 
    -- predecessors 52 55 
    -- successors 56 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_48 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(52);
      predecessors(1) <= cp_elements(55);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(48)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(48),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => array_obj_ref_606_index_sum_1_req_0); -- 
    -- CP-element group 49 transition  output  bypass 
    -- predecessors 37 
    -- successors 50 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_604_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_604_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_604_completed_
      -- 
    cp_elements(49) <= cp_elements(37);
    index_resize_req_1467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => array_obj_ref_606_index_0_resize_req_0); -- 
    -- CP-element group 50 transition  input  output  no-bypass 
    -- predecessors 49 
    -- successors 51 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_0_resize_ack_0, ack => cp_elements(50)); -- 
    scale_rr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => array_obj_ref_606_index_0_scale_req_0); -- 
    -- CP-element group 51 transition  input  output  no-bypass 
    -- predecessors 50 
    -- successors 52 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_0/scale_cr
      -- 
    scale_ra_1473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_0_scale_ack_0, ack => cp_elements(51)); -- 
    scale_cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => array_obj_ref_606_index_0_scale_req_1); -- 
    -- CP-element group 52 transition  input  no-bypass 
    -- predecessors 51 
    -- successors 48 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_0/scale_ca
      -- 
    scale_ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_0_scale_ack_1, ack => cp_elements(52)); -- 
    -- CP-element group 53 transition  output  bypass 
    -- predecessors 39 
    -- successors 54 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_605_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_605_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_605_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_1/index_resize_req
      -- 
    cp_elements(53) <= cp_elements(39);
    index_resize_req_1484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => array_obj_ref_606_index_1_resize_req_0); -- 
    -- CP-element group 54 transition  input  output  no-bypass 
    -- predecessors 53 
    -- successors 55 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_1485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_1_resize_ack_0, ack => cp_elements(54)); -- 
    scale_rename_req_1489_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => array_obj_ref_606_index_1_rename_req_0); -- 
    -- CP-element group 55 transition  input  no-bypass 
    -- predecessors 54 
    -- successors 48 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_1490_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_1_rename_ack_0, ack => cp_elements(55)); -- 
    -- CP-element group 56 transition  input  output  no-bypass 
    -- predecessors 48 
    -- successors 57 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_1495_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_sum_1_ack_0, ack => cp_elements(56)); -- 
    partial_sum_1_cr_1496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => array_obj_ref_606_index_sum_1_req_1); -- 
    -- CP-element group 57 transition  input  output  no-bypass 
    -- predecessors 56 
    -- successors 58 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/final_index_req
      -- 
    partial_sum_1_ca_1497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_sum_1_ack_1, ack => cp_elements(57)); -- 
    final_index_req_1498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => array_obj_ref_606_offset_inst_req_0); -- 
    -- CP-element group 58 transition  input  output  no-bypass 
    -- predecessors 57 
    -- successors 59 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_add_indices/$exit
      -- 
    final_index_ack_1499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_offset_inst_ack_0, ack => cp_elements(58)); -- 
    sum_rename_req_1503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => array_obj_ref_606_root_address_inst_req_0); -- 
    -- CP-element group 59 transition  input  no-bypass 
    -- predecessors 58 
    -- successors 46 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_606_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_root_address_inst_ack_0, ack => cp_elements(59)); -- 
    -- CP-element group 60 transition  output  bypass 
    -- predecessors 46 
    -- successors 61 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_607_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_607_complete/final_reg_req
      -- 
    cp_elements(60) <= cp_elements(46);
    final_reg_req_1508_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => addr_of_607_final_reg_req_0); -- 
    -- CP-element group 61 transition  input  no-bypass 
    -- predecessors 60 
    -- successors 47 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_607_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_607_complete/final_reg_ack
      -- 
    final_reg_ack_1509_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_607_final_reg_ack_0, ack => cp_elements(61)); -- 
    -- CP-element group 62 join  fork  transition  no-bypass 
    -- predecessors 64 66 
    -- successors 63 67 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_active_
      -- 
    cpelement_group_62 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(64);
      predecessors(1) <= cp_elements(66);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(62)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(62),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 63 join  fork  transition  no-bypass 
    -- predecessors 62 68 
    -- successors 77 135 210 278 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_614_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_614_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_614_completed_
      -- 
    cpelement_group_63 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(62);
      predecessors(1) <= cp_elements(68);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(63)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(63),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 64 fork  transition  bypass 
    -- predecessors 39 
    -- successors 62 65 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_610_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_610_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_610_completed_
      -- 
    cp_elements(64) <= cp_elements(39);
    -- CP-element group 65 transition  output  bypass 
    -- predecessors 64 
    -- successors 66 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Sample/rr
      -- 
    cp_elements(65) <= cp_elements(64);
    rr_1522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => binary_613_inst_req_0); -- 
    -- CP-element group 66 transition  input  no-bypass 
    -- predecessors 65 
    -- successors 62 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Sample/ra
      -- 
    ra_1523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_613_inst_ack_0, ack => cp_elements(66)); -- 
    -- CP-element group 67 transition  output  bypass 
    -- predecessors 62 
    -- successors 68 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Update/cr
      -- 
    cp_elements(67) <= cp_elements(62);
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => binary_613_inst_req_1); -- 
    -- CP-element group 68 transition  input  no-bypass 
    -- predecessors 67 
    -- successors 63 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_613_complete_Update/$exit
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_613_inst_ack_1, ack => cp_elements(68)); -- 
    -- CP-element group 69 transition  bypass 
    -- predecessors 37 
    -- successors 70 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_619_trigger_
      -- 
    cp_elements(69) <= cp_elements(37);
    -- CP-element group 70 join  fork  transition  bypass 
    -- predecessors 69 83 
    -- successors 71 84 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_619_active_
      -- 
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(69);
      predecessors(1) <= cp_elements(83);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(70)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 71 join  transition  no-bypass 
    -- predecessors 70 85 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_620_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_620_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_620_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_619_completed_
      -- 
    cpelement_group_71 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(70);
      predecessors(1) <= cp_elements(85);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(71)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(71),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 72 join  transition  output  bypass 
    -- predecessors 76 79 
    -- successors 80 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(76);
      predecessors(1) <= cp_elements(79);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(72)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_618_index_sum_1_req_0); -- 
    -- CP-element group 73 transition  output  bypass 
    -- predecessors 37 
    -- successors 74 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_616_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_616_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_616_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_computed_0
      -- 
    cp_elements(73) <= cp_elements(37);
    index_resize_req_1546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => array_obj_ref_618_index_0_resize_req_0); -- 
    -- CP-element group 74 transition  input  output  no-bypass 
    -- predecessors 73 
    -- successors 75 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_index_0_resize_ack_0, ack => cp_elements(74)); -- 
    scale_rr_1551_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => array_obj_ref_618_index_0_scale_req_0); -- 
    -- CP-element group 75 transition  input  output  no-bypass 
    -- predecessors 74 
    -- successors 76 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_0/scale_ra
      -- 
    scale_ra_1552_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_index_0_scale_ack_0, ack => cp_elements(75)); -- 
    scale_cr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => array_obj_ref_618_index_0_scale_req_1); -- 
    -- CP-element group 76 transition  input  no-bypass 
    -- predecessors 75 
    -- successors 72 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_0/$exit
      -- 
    scale_ca_1554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_index_0_scale_ack_1, ack => cp_elements(76)); -- 
    -- CP-element group 77 transition  output  bypass 
    -- predecessors 63 
    -- successors 78 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_617_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_617_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_617_completed_
      -- 
    cp_elements(77) <= cp_elements(63);
    index_resize_req_1563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => array_obj_ref_618_index_1_resize_req_0); -- 
    -- CP-element group 78 transition  input  output  no-bypass 
    -- predecessors 77 
    -- successors 79 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_1/$entry
      -- 
    index_resize_ack_1564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_index_1_resize_ack_0, ack => cp_elements(78)); -- 
    scale_rename_req_1568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => array_obj_ref_618_index_1_rename_req_0); -- 
    -- CP-element group 79 transition  input  no-bypass 
    -- predecessors 78 
    -- successors 72 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_1569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_index_1_rename_ack_0, ack => cp_elements(79)); -- 
    -- CP-element group 80 transition  input  output  no-bypass 
    -- predecessors 72 
    -- successors 81 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_1574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_index_sum_1_ack_0, ack => cp_elements(80)); -- 
    partial_sum_1_cr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => array_obj_ref_618_index_sum_1_req_1); -- 
    -- CP-element group 81 transition  input  output  no-bypass 
    -- predecessors 80 
    -- successors 82 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_1576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_index_sum_1_ack_1, ack => cp_elements(81)); -- 
    final_index_req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => array_obj_ref_618_offset_inst_req_0); -- 
    -- CP-element group 82 transition  input  output  no-bypass 
    -- predecessors 81 
    -- successors 83 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_add_indices/final_index_ack
      -- 
    final_index_ack_1578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_offset_inst_ack_0, ack => cp_elements(82)); -- 
    sum_rename_req_1582_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => array_obj_ref_618_root_address_inst_req_0); -- 
    -- CP-element group 83 transition  input  no-bypass 
    -- predecessors 82 
    -- successors 70 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_618_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1583_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_618_root_address_inst_ack_0, ack => cp_elements(83)); -- 
    -- CP-element group 84 transition  output  bypass 
    -- predecessors 70 
    -- successors 85 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_619_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_619_complete/$entry
      -- 
    cp_elements(84) <= cp_elements(70);
    final_reg_req_1587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => addr_of_619_final_reg_req_0); -- 
    -- CP-element group 85 transition  input  no-bypass 
    -- predecessors 84 
    -- successors 71 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_619_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_619_complete/final_reg_ack
      -- 
    final_reg_ack_1588_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_619_final_reg_ack_0, ack => cp_elements(85)); -- 
    -- CP-element group 86 join  fork  transition  no-bypass 
    -- predecessors 88 90 
    -- successors 87 91 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_active_
      -- 
    cpelement_group_86 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(88);
      predecessors(1) <= cp_elements(90);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(86)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(86),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 87 join  fork  transition  no-bypass 
    -- predecessors 86 92 
    -- successors 101 152 227 295 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_626_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_626_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_626_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_completed_
      -- 
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(86);
      predecessors(1) <= cp_elements(92);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(87)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 88 fork  transition  bypass 
    -- predecessors 39 
    -- successors 86 89 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_622_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_622_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_622_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_trigger_
      -- 
    cp_elements(88) <= cp_elements(39);
    -- CP-element group 89 transition  output  bypass 
    -- predecessors 88 
    -- successors 90 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Sample/$entry
      -- 
    cp_elements(89) <= cp_elements(88);
    rr_1601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => binary_625_inst_req_0); -- 
    -- CP-element group 90 transition  input  no-bypass 
    -- predecessors 89 
    -- successors 86 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Sample/ra
      -- 
    ra_1602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_625_inst_ack_0, ack => cp_elements(90)); -- 
    -- CP-element group 91 transition  output  bypass 
    -- predecessors 86 
    -- successors 92 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Update/cr
      -- 
    cp_elements(91) <= cp_elements(86);
    cr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => binary_625_inst_req_1); -- 
    -- CP-element group 92 transition  input  no-bypass 
    -- predecessors 91 
    -- successors 87 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_625_complete_Update/$exit
      -- 
    ca_1607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_625_inst_ack_1, ack => cp_elements(92)); -- 
    -- CP-element group 93 transition  bypass 
    -- predecessors 37 
    -- successors 94 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_631_trigger_
      -- 
    cp_elements(93) <= cp_elements(37);
    -- CP-element group 94 join  fork  transition  bypass 
    -- predecessors 93 107 
    -- successors 95 108 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_631_active_
      -- 
    cpelement_group_94 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(93);
      predecessors(1) <= cp_elements(107);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(94)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(94),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 95 join  transition  no-bypass 
    -- predecessors 94 109 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_631_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_632_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_632_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_632_trigger_
      -- 
    cpelement_group_95 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(94);
      predecessors(1) <= cp_elements(109);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(95)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(95),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 96 join  transition  output  bypass 
    -- predecessors 100 103 
    -- successors 104 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_indices_scaled
      -- 
    cpelement_group_96 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(100);
      predecessors(1) <= cp_elements(103);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(96)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(96),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1652_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => array_obj_ref_630_index_sum_1_req_0); -- 
    -- CP-element group 97 transition  output  bypass 
    -- predecessors 37 
    -- successors 98 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_628_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_628_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_628_trigger_
      -- 
    cp_elements(97) <= cp_elements(37);
    index_resize_req_1625_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => array_obj_ref_630_index_0_resize_req_0); -- 
    -- CP-element group 98 transition  input  output  no-bypass 
    -- predecessors 97 
    -- successors 99 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_0/scale_rr
      -- 
    index_resize_ack_1626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_index_0_resize_ack_0, ack => cp_elements(98)); -- 
    scale_rr_1630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => array_obj_ref_630_index_0_scale_req_0); -- 
    -- CP-element group 99 transition  input  output  no-bypass 
    -- predecessors 98 
    -- successors 100 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_0/scale_ra
      -- 
    scale_ra_1631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_index_0_scale_ack_0, ack => cp_elements(99)); -- 
    scale_cr_1632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => array_obj_ref_630_index_0_scale_req_1); -- 
    -- CP-element group 100 transition  input  no-bypass 
    -- predecessors 99 
    -- successors 96 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_0/$exit
      -- 
    scale_ca_1633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_index_0_scale_ack_1, ack => cp_elements(100)); -- 
    -- CP-element group 101 transition  output  bypass 
    -- predecessors 87 
    -- successors 102 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_629_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_629_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_629_completed_
      -- 
    cp_elements(101) <= cp_elements(87);
    index_resize_req_1642_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => array_obj_ref_630_index_1_resize_req_0); -- 
    -- CP-element group 102 transition  input  output  no-bypass 
    -- predecessors 101 
    -- successors 103 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_resize_1/index_resize_ack
      -- 
    index_resize_ack_1643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_index_1_resize_ack_0, ack => cp_elements(102)); -- 
    scale_rename_req_1647_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => array_obj_ref_630_index_1_rename_req_0); -- 
    -- CP-element group 103 transition  input  no-bypass 
    -- predecessors 102 
    -- successors 96 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_index_scale_1/$exit
      -- 
    scale_rename_ack_1648_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_index_1_rename_ack_0, ack => cp_elements(103)); -- 
    -- CP-element group 104 transition  input  output  no-bypass 
    -- predecessors 96 
    -- successors 105 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_1653_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_index_sum_1_ack_0, ack => cp_elements(104)); -- 
    partial_sum_1_cr_1654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => array_obj_ref_630_index_sum_1_req_1); -- 
    -- CP-element group 105 transition  input  output  no-bypass 
    -- predecessors 104 
    -- successors 106 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/final_index_req
      -- 
    partial_sum_1_ca_1655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_index_sum_1_ack_1, ack => cp_elements(105)); -- 
    final_index_req_1656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => array_obj_ref_630_offset_inst_req_0); -- 
    -- CP-element group 106 transition  input  output  no-bypass 
    -- predecessors 105 
    -- successors 107 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_offset_calculated
      -- 
    final_index_ack_1657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_offset_inst_ack_0, ack => cp_elements(106)); -- 
    sum_rename_req_1661_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => array_obj_ref_630_root_address_inst_req_0); -- 
    -- CP-element group 107 transition  input  no-bypass 
    -- predecessors 106 
    -- successors 94 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_630_root_address_calculated
      -- 
    sum_rename_ack_1662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_630_root_address_inst_ack_0, ack => cp_elements(107)); -- 
    -- CP-element group 108 transition  output  bypass 
    -- predecessors 94 
    -- successors 109 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_631_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_631_complete/final_reg_req
      -- 
    cp_elements(108) <= cp_elements(94);
    final_reg_req_1666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => addr_of_631_final_reg_req_0); -- 
    -- CP-element group 109 transition  input  no-bypass 
    -- predecessors 108 
    -- successors 95 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_631_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_631_complete/final_reg_ack
      -- 
    final_reg_ack_1667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_631_final_reg_ack_0, ack => cp_elements(109)); -- 
    -- CP-element group 110 transition  bypass 
    -- predecessors 37 
    -- successors 111 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_637_trigger_
      -- 
    cp_elements(110) <= cp_elements(37);
    -- CP-element group 111 join  fork  transition  bypass 
    -- predecessors 110 124 
    -- successors 112 125 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_637_active_
      -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(110);
      predecessors(1) <= cp_elements(124);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(111)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 112 join  transition  no-bypass 
    -- predecessors 111 126 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_637_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_638_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_638_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_638_active_
      -- 
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(111);
      predecessors(1) <= cp_elements(126);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(112)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 113 join  transition  output  bypass 
    -- predecessors 117 120 
    -- successors 121 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_113 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(117);
      predecessors(1) <= cp_elements(120);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(113)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => array_obj_ref_636_index_sum_1_req_0); -- 
    -- CP-element group 114 transition  output  bypass 
    -- predecessors 37 
    -- successors 115 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_634_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_634_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_634_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_0/index_resize_req
      -- 
    cp_elements(114) <= cp_elements(37);
    index_resize_req_1685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => array_obj_ref_636_index_0_resize_req_0); -- 
    -- CP-element group 115 transition  input  output  no-bypass 
    -- predecessors 114 
    -- successors 116 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_0/scale_rr
      -- 
    index_resize_ack_1686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_index_0_resize_ack_0, ack => cp_elements(115)); -- 
    scale_rr_1690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_636_index_0_scale_req_0); -- 
    -- CP-element group 116 transition  input  output  no-bypass 
    -- predecessors 115 
    -- successors 117 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_0/scale_cr
      -- 
    scale_ra_1691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_index_0_scale_ack_0, ack => cp_elements(116)); -- 
    scale_cr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_636_index_0_scale_req_1); -- 
    -- CP-element group 117 transition  input  no-bypass 
    -- predecessors 116 
    -- successors 113 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_0/scale_ca
      -- 
    scale_ca_1693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_index_0_scale_ack_1, ack => cp_elements(117)); -- 
    -- CP-element group 118 transition  output  bypass 
    -- predecessors 39 
    -- successors 119 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_635_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_635_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_635_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_1/index_resize_req
      -- 
    cp_elements(118) <= cp_elements(39);
    index_resize_req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_636_index_1_resize_req_0); -- 
    -- CP-element group 119 transition  input  output  no-bypass 
    -- predecessors 118 
    -- successors 120 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_1703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_index_1_resize_ack_0, ack => cp_elements(119)); -- 
    scale_rename_req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => array_obj_ref_636_index_1_rename_req_0); -- 
    -- CP-element group 120 transition  input  no-bypass 
    -- predecessors 119 
    -- successors 113 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_1708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_index_1_rename_ack_0, ack => cp_elements(120)); -- 
    -- CP-element group 121 transition  input  output  no-bypass 
    -- predecessors 113 
    -- successors 122 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_1713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_index_sum_1_ack_0, ack => cp_elements(121)); -- 
    partial_sum_1_cr_1714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => array_obj_ref_636_index_sum_1_req_1); -- 
    -- CP-element group 122 transition  input  output  no-bypass 
    -- predecessors 121 
    -- successors 123 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/final_index_req
      -- 
    partial_sum_1_ca_1715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_index_sum_1_ack_1, ack => cp_elements(122)); -- 
    final_index_req_1716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => array_obj_ref_636_offset_inst_req_0); -- 
    -- CP-element group 123 transition  input  output  no-bypass 
    -- predecessors 122 
    -- successors 124 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_1717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_offset_inst_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_1721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => array_obj_ref_636_root_address_inst_req_0); -- 
    -- CP-element group 124 transition  input  no-bypass 
    -- predecessors 123 
    -- successors 111 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_636_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_636_root_address_inst_ack_0, ack => cp_elements(124)); -- 
    -- CP-element group 125 transition  output  bypass 
    -- predecessors 111 
    -- successors 126 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_637_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_637_complete/final_reg_req
      -- 
    cp_elements(125) <= cp_elements(111);
    final_reg_req_1726_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => addr_of_637_final_reg_req_0); -- 
    -- CP-element group 126 transition  input  no-bypass 
    -- predecessors 125 
    -- successors 112 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_637_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_637_complete/final_reg_ack
      -- 
    final_reg_ack_1727_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_637_final_reg_ack_0, ack => cp_elements(126)); -- 
    -- CP-element group 127 transition  bypass 
    -- predecessors 37 
    -- successors 128 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_643_trigger_
      -- 
    cp_elements(127) <= cp_elements(37);
    -- CP-element group 128 join  fork  transition  bypass 
    -- predecessors 127 141 
    -- successors 129 142 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_643_active_
      -- 
    cpelement_group_128 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(127);
      predecessors(1) <= cp_elements(141);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(128)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(128),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 129 join  transition  no-bypass 
    -- predecessors 128 143 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_644_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_644_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_644_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_643_completed_
      -- 
    cpelement_group_129 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(128);
      predecessors(1) <= cp_elements(143);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(129)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(129),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 130 join  transition  output  bypass 
    -- predecessors 134 137 
    -- successors 138 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_130 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(134);
      predecessors(1) <= cp_elements(137);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(130)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => array_obj_ref_642_index_sum_1_req_0); -- 
    -- CP-element group 131 transition  output  bypass 
    -- predecessors 37 
    -- successors 132 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_640_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_640_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_640_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_0/index_resize_req
      -- 
    cp_elements(131) <= cp_elements(37);
    index_resize_req_1745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => array_obj_ref_642_index_0_resize_req_0); -- 
    -- CP-element group 132 transition  input  output  no-bypass 
    -- predecessors 131 
    -- successors 133 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_0/scale_rr
      -- 
    index_resize_ack_1746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_index_0_resize_ack_0, ack => cp_elements(132)); -- 
    scale_rr_1750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => array_obj_ref_642_index_0_scale_req_0); -- 
    -- CP-element group 133 transition  input  output  no-bypass 
    -- predecessors 132 
    -- successors 134 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_0/scale_cr
      -- 
    scale_ra_1751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_index_0_scale_ack_0, ack => cp_elements(133)); -- 
    scale_cr_1752_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(133), ack => array_obj_ref_642_index_0_scale_req_1); -- 
    -- CP-element group 134 transition  input  no-bypass 
    -- predecessors 133 
    -- successors 130 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_0/scale_ca
      -- 
    scale_ca_1753_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_index_0_scale_ack_1, ack => cp_elements(134)); -- 
    -- CP-element group 135 transition  output  bypass 
    -- predecessors 63 
    -- successors 136 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_641_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_641_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_641_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_1/index_resize_req
      -- 
    cp_elements(135) <= cp_elements(63);
    index_resize_req_1762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => array_obj_ref_642_index_1_resize_req_0); -- 
    -- CP-element group 136 transition  input  output  no-bypass 
    -- predecessors 135 
    -- successors 137 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_1763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_index_1_resize_ack_0, ack => cp_elements(136)); -- 
    scale_rename_req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => array_obj_ref_642_index_1_rename_req_0); -- 
    -- CP-element group 137 transition  input  no-bypass 
    -- predecessors 136 
    -- successors 130 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_index_1_rename_ack_0, ack => cp_elements(137)); -- 
    -- CP-element group 138 transition  input  output  no-bypass 
    -- predecessors 130 
    -- successors 139 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_1773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_index_sum_1_ack_0, ack => cp_elements(138)); -- 
    partial_sum_1_cr_1774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => array_obj_ref_642_index_sum_1_req_1); -- 
    -- CP-element group 139 transition  input  output  no-bypass 
    -- predecessors 138 
    -- successors 140 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/final_index_req
      -- 
    partial_sum_1_ca_1775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_index_sum_1_ack_1, ack => cp_elements(139)); -- 
    final_index_req_1776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => array_obj_ref_642_offset_inst_req_0); -- 
    -- CP-element group 140 transition  input  output  no-bypass 
    -- predecessors 139 
    -- successors 141 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_1777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_offset_inst_ack_0, ack => cp_elements(140)); -- 
    sum_rename_req_1781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => array_obj_ref_642_root_address_inst_req_0); -- 
    -- CP-element group 141 transition  input  no-bypass 
    -- predecessors 140 
    -- successors 128 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_642_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_642_root_address_inst_ack_0, ack => cp_elements(141)); -- 
    -- CP-element group 142 transition  output  bypass 
    -- predecessors 128 
    -- successors 143 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_643_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_643_complete/final_reg_req
      -- 
    cp_elements(142) <= cp_elements(128);
    final_reg_req_1786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => addr_of_643_final_reg_req_0); -- 
    -- CP-element group 143 transition  input  no-bypass 
    -- predecessors 142 
    -- successors 129 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_643_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_643_complete/final_reg_ack
      -- 
    final_reg_ack_1787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_643_final_reg_ack_0, ack => cp_elements(143)); -- 
    -- CP-element group 144 transition  bypass 
    -- predecessors 37 
    -- successors 145 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_649_trigger_
      -- 
    cp_elements(144) <= cp_elements(37);
    -- CP-element group 145 join  fork  transition  bypass 
    -- predecessors 144 158 
    -- successors 146 159 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_649_active_
      -- 
    cpelement_group_145 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(144);
      predecessors(1) <= cp_elements(158);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(145)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(145),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 146 join  transition  no-bypass 
    -- predecessors 145 160 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_650_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_650_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_650_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_649_completed_
      -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(145);
      predecessors(1) <= cp_elements(160);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(146)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 147 join  transition  output  bypass 
    -- predecessors 151 154 
    -- successors 155 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_147 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(151);
      predecessors(1) <= cp_elements(154);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(147)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => array_obj_ref_648_index_sum_1_req_0); -- 
    -- CP-element group 148 transition  output  bypass 
    -- predecessors 37 
    -- successors 149 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_646_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_646_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_646_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_0/index_resize_req
      -- 
    cp_elements(148) <= cp_elements(37);
    index_resize_req_1805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => array_obj_ref_648_index_0_resize_req_0); -- 
    -- CP-element group 149 transition  input  output  no-bypass 
    -- predecessors 148 
    -- successors 150 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_0/scale_rr
      -- 
    index_resize_ack_1806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_index_0_resize_ack_0, ack => cp_elements(149)); -- 
    scale_rr_1810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => array_obj_ref_648_index_0_scale_req_0); -- 
    -- CP-element group 150 transition  input  output  no-bypass 
    -- predecessors 149 
    -- successors 151 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_0/scale_cr
      -- 
    scale_ra_1811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_index_0_scale_ack_0, ack => cp_elements(150)); -- 
    scale_cr_1812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(150), ack => array_obj_ref_648_index_0_scale_req_1); -- 
    -- CP-element group 151 transition  input  no-bypass 
    -- predecessors 150 
    -- successors 147 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_0/scale_ca
      -- 
    scale_ca_1813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_index_0_scale_ack_1, ack => cp_elements(151)); -- 
    -- CP-element group 152 transition  output  bypass 
    -- predecessors 87 
    -- successors 153 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_647_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_647_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_647_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_1/index_resize_req
      -- 
    cp_elements(152) <= cp_elements(87);
    index_resize_req_1822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(152), ack => array_obj_ref_648_index_1_resize_req_0); -- 
    -- CP-element group 153 transition  input  output  no-bypass 
    -- predecessors 152 
    -- successors 154 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_1823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_index_1_resize_ack_0, ack => cp_elements(153)); -- 
    scale_rename_req_1827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => array_obj_ref_648_index_1_rename_req_0); -- 
    -- CP-element group 154 transition  input  no-bypass 
    -- predecessors 153 
    -- successors 147 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_1828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_index_1_rename_ack_0, ack => cp_elements(154)); -- 
    -- CP-element group 155 transition  input  output  no-bypass 
    -- predecessors 147 
    -- successors 156 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_1833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_index_sum_1_ack_0, ack => cp_elements(155)); -- 
    partial_sum_1_cr_1834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => array_obj_ref_648_index_sum_1_req_1); -- 
    -- CP-element group 156 transition  input  output  no-bypass 
    -- predecessors 155 
    -- successors 157 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/final_index_req
      -- 
    partial_sum_1_ca_1835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_index_sum_1_ack_1, ack => cp_elements(156)); -- 
    final_index_req_1836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(156), ack => array_obj_ref_648_offset_inst_req_0); -- 
    -- CP-element group 157 transition  input  output  no-bypass 
    -- predecessors 156 
    -- successors 158 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_1837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_offset_inst_ack_0, ack => cp_elements(157)); -- 
    sum_rename_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => array_obj_ref_648_root_address_inst_req_0); -- 
    -- CP-element group 158 transition  input  no-bypass 
    -- predecessors 157 
    -- successors 145 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_648_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_648_root_address_inst_ack_0, ack => cp_elements(158)); -- 
    -- CP-element group 159 transition  output  bypass 
    -- predecessors 145 
    -- successors 160 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_649_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_649_complete/final_reg_req
      -- 
    cp_elements(159) <= cp_elements(145);
    final_reg_req_1846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(159), ack => addr_of_649_final_reg_req_0); -- 
    -- CP-element group 160 transition  input  no-bypass 
    -- predecessors 159 
    -- successors 146 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_649_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_649_complete/final_reg_ack
      -- 
    final_reg_ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_649_final_reg_ack_0, ack => cp_elements(160)); -- 
    -- CP-element group 161 join  fork  transition  no-bypass 
    -- predecessors 163 165 
    -- successors 162 166 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_active_
      -- 
    cpelement_group_161 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(163);
      predecessors(1) <= cp_elements(165);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(161)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(161),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 162 join  fork  transition  no-bypass 
    -- predecessors 161 167 
    -- successors 176 244 312 329 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_656_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_656_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_656_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_completed_
      -- 
    cpelement_group_162 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(161);
      predecessors(1) <= cp_elements(167);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(162)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(162),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 163 fork  transition  bypass 
    -- predecessors 39 
    -- successors 161 164 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_652_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_652_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_652_completed_
      -- 
    cp_elements(163) <= cp_elements(39);
    -- CP-element group 164 transition  output  bypass 
    -- predecessors 163 
    -- successors 165 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Sample/rr
      -- 
    cp_elements(164) <= cp_elements(163);
    rr_1860_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => binary_655_inst_req_0); -- 
    -- CP-element group 165 transition  input  no-bypass 
    -- predecessors 164 
    -- successors 161 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Sample/ra
      -- 
    ra_1861_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_655_inst_ack_0, ack => cp_elements(165)); -- 
    -- CP-element group 166 transition  output  bypass 
    -- predecessors 161 
    -- successors 167 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Update/cr
      -- 
    cp_elements(166) <= cp_elements(161);
    cr_1865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => binary_655_inst_req_1); -- 
    -- CP-element group 167 transition  input  no-bypass 
    -- predecessors 166 
    -- successors 162 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_655_complete_Update/ca
      -- 
    ca_1866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_655_inst_ack_1, ack => cp_elements(167)); -- 
    -- CP-element group 168 transition  bypass 
    -- predecessors 37 
    -- successors 169 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_661_trigger_
      -- 
    cp_elements(168) <= cp_elements(37);
    -- CP-element group 169 join  fork  transition  bypass 
    -- predecessors 168 182 
    -- successors 170 183 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_661_active_
      -- 
    cpelement_group_169 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(168);
      predecessors(1) <= cp_elements(182);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(169)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(169),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 170 join  transition  no-bypass 
    -- predecessors 169 184 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_662_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_662_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_662_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_661_completed_
      -- 
    cpelement_group_170 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(169);
      predecessors(1) <= cp_elements(184);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(170)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(170),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 171 join  transition  output  bypass 
    -- predecessors 175 178 
    -- successors 179 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_171 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(175);
      predecessors(1) <= cp_elements(178);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(171)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(171),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1911_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => array_obj_ref_660_index_sum_1_req_0); -- 
    -- CP-element group 172 transition  output  bypass 
    -- predecessors 37 
    -- successors 173 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_658_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_658_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_658_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_0/index_resize_req
      -- 
    cp_elements(172) <= cp_elements(37);
    index_resize_req_1884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(172), ack => array_obj_ref_660_index_0_resize_req_0); -- 
    -- CP-element group 173 transition  input  output  no-bypass 
    -- predecessors 172 
    -- successors 174 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_0/scale_rr
      -- 
    index_resize_ack_1885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_0_resize_ack_0, ack => cp_elements(173)); -- 
    scale_rr_1889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => array_obj_ref_660_index_0_scale_req_0); -- 
    -- CP-element group 174 transition  input  output  no-bypass 
    -- predecessors 173 
    -- successors 175 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_0/scale_cr
      -- 
    scale_ra_1890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_0_scale_ack_0, ack => cp_elements(174)); -- 
    scale_cr_1891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(174), ack => array_obj_ref_660_index_0_scale_req_1); -- 
    -- CP-element group 175 transition  input  no-bypass 
    -- predecessors 174 
    -- successors 171 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_0/scale_ca
      -- 
    scale_ca_1892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_0_scale_ack_1, ack => cp_elements(175)); -- 
    -- CP-element group 176 transition  output  bypass 
    -- predecessors 162 
    -- successors 177 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_659_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_659_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_659_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_1/index_resize_req
      -- 
    cp_elements(176) <= cp_elements(162);
    index_resize_req_1901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => array_obj_ref_660_index_1_resize_req_0); -- 
    -- CP-element group 177 transition  input  output  no-bypass 
    -- predecessors 176 
    -- successors 178 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_1902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_1_resize_ack_0, ack => cp_elements(177)); -- 
    scale_rename_req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => array_obj_ref_660_index_1_rename_req_0); -- 
    -- CP-element group 178 transition  input  no-bypass 
    -- predecessors 177 
    -- successors 171 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_1_rename_ack_0, ack => cp_elements(178)); -- 
    -- CP-element group 179 transition  input  output  no-bypass 
    -- predecessors 171 
    -- successors 180 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_1912_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_sum_1_ack_0, ack => cp_elements(179)); -- 
    partial_sum_1_cr_1913_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => array_obj_ref_660_index_sum_1_req_1); -- 
    -- CP-element group 180 transition  input  output  no-bypass 
    -- predecessors 179 
    -- successors 181 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/final_index_req
      -- 
    partial_sum_1_ca_1914_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_sum_1_ack_1, ack => cp_elements(180)); -- 
    final_index_req_1915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => array_obj_ref_660_offset_inst_req_0); -- 
    -- CP-element group 181 transition  input  output  no-bypass 
    -- predecessors 180 
    -- successors 182 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_1916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_offset_inst_ack_0, ack => cp_elements(181)); -- 
    sum_rename_req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => array_obj_ref_660_root_address_inst_req_0); -- 
    -- CP-element group 182 transition  input  no-bypass 
    -- predecessors 181 
    -- successors 169 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_660_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_root_address_inst_ack_0, ack => cp_elements(182)); -- 
    -- CP-element group 183 transition  output  bypass 
    -- predecessors 169 
    -- successors 184 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_661_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_661_complete/final_reg_req
      -- 
    cp_elements(183) <= cp_elements(169);
    final_reg_req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => addr_of_661_final_reg_req_0); -- 
    -- CP-element group 184 transition  input  no-bypass 
    -- predecessors 183 
    -- successors 170 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_661_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_661_complete/final_reg_ack
      -- 
    final_reg_ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_661_final_reg_ack_0, ack => cp_elements(184)); -- 
    -- CP-element group 185 transition  bypass 
    -- predecessors 37 
    -- successors 186 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_667_trigger_
      -- 
    cp_elements(185) <= cp_elements(37);
    -- CP-element group 186 join  fork  transition  bypass 
    -- predecessors 185 199 
    -- successors 187 200 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_667_active_
      -- 
    cpelement_group_186 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(185);
      predecessors(1) <= cp_elements(199);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(186)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(186),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 187 join  transition  no-bypass 
    -- predecessors 186 201 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_668_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_668_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_668_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_667_completed_
      -- 
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(186);
      predecessors(1) <= cp_elements(201);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(187)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 188 join  transition  output  bypass 
    -- predecessors 192 195 
    -- successors 196 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_188 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(192);
      predecessors(1) <= cp_elements(195);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(188)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(188),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_1971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => array_obj_ref_666_index_sum_1_req_0); -- 
    -- CP-element group 189 transition  output  bypass 
    -- predecessors 37 
    -- successors 190 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_664_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_664_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_664_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_0/index_resize_req
      -- 
    cp_elements(189) <= cp_elements(37);
    index_resize_req_1944_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => array_obj_ref_666_index_0_resize_req_0); -- 
    -- CP-element group 190 transition  input  output  no-bypass 
    -- predecessors 189 
    -- successors 191 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_0/scale_rr
      -- 
    index_resize_ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_index_0_resize_ack_0, ack => cp_elements(190)); -- 
    scale_rr_1949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => array_obj_ref_666_index_0_scale_req_0); -- 
    -- CP-element group 191 transition  input  output  no-bypass 
    -- predecessors 190 
    -- successors 192 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_0/scale_cr
      -- 
    scale_ra_1950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_index_0_scale_ack_0, ack => cp_elements(191)); -- 
    scale_cr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(191), ack => array_obj_ref_666_index_0_scale_req_1); -- 
    -- CP-element group 192 transition  input  no-bypass 
    -- predecessors 191 
    -- successors 188 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_0/scale_ca
      -- 
    scale_ca_1952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_index_0_scale_ack_1, ack => cp_elements(192)); -- 
    -- CP-element group 193 transition  output  bypass 
    -- predecessors 39 
    -- successors 194 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_665_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_665_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_665_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_1/index_resize_req
      -- 
    cp_elements(193) <= cp_elements(39);
    index_resize_req_1961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => array_obj_ref_666_index_1_resize_req_0); -- 
    -- CP-element group 194 transition  input  output  no-bypass 
    -- predecessors 193 
    -- successors 195 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_1962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_index_1_resize_ack_0, ack => cp_elements(194)); -- 
    scale_rename_req_1966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => array_obj_ref_666_index_1_rename_req_0); -- 
    -- CP-element group 195 transition  input  no-bypass 
    -- predecessors 194 
    -- successors 188 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_1967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_index_1_rename_ack_0, ack => cp_elements(195)); -- 
    -- CP-element group 196 transition  input  output  no-bypass 
    -- predecessors 188 
    -- successors 197 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_1972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_index_sum_1_ack_0, ack => cp_elements(196)); -- 
    partial_sum_1_cr_1973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => array_obj_ref_666_index_sum_1_req_1); -- 
    -- CP-element group 197 transition  input  output  no-bypass 
    -- predecessors 196 
    -- successors 198 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/final_index_req
      -- 
    partial_sum_1_ca_1974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_index_sum_1_ack_1, ack => cp_elements(197)); -- 
    final_index_req_1975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => array_obj_ref_666_offset_inst_req_0); -- 
    -- CP-element group 198 transition  input  output  no-bypass 
    -- predecessors 197 
    -- successors 199 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_offset_inst_ack_0, ack => cp_elements(198)); -- 
    sum_rename_req_1980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => array_obj_ref_666_root_address_inst_req_0); -- 
    -- CP-element group 199 transition  input  no-bypass 
    -- predecessors 198 
    -- successors 186 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_666_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_666_root_address_inst_ack_0, ack => cp_elements(199)); -- 
    -- CP-element group 200 transition  output  bypass 
    -- predecessors 186 
    -- successors 201 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_667_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_667_complete/final_reg_req
      -- 
    cp_elements(200) <= cp_elements(186);
    final_reg_req_1985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => addr_of_667_final_reg_req_0); -- 
    -- CP-element group 201 transition  input  no-bypass 
    -- predecessors 200 
    -- successors 187 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_667_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_667_complete/final_reg_ack
      -- 
    final_reg_ack_1986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_667_final_reg_ack_0, ack => cp_elements(201)); -- 
    -- CP-element group 202 transition  bypass 
    -- predecessors 37 
    -- successors 203 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_673_trigger_
      -- 
    cp_elements(202) <= cp_elements(37);
    -- CP-element group 203 join  fork  transition  bypass 
    -- predecessors 202 216 
    -- successors 204 217 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_673_active_
      -- 
    cpelement_group_203 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(202);
      predecessors(1) <= cp_elements(216);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(203)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(203),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 204 join  transition  no-bypass 
    -- predecessors 203 218 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_673_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_674_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_674_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_674_completed_
      -- 
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(203);
      predecessors(1) <= cp_elements(218);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(204)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 205 join  transition  output  bypass 
    -- predecessors 209 212 
    -- successors 213 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_indices_scaled
      -- 
    cpelement_group_205 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(209);
      predecessors(1) <= cp_elements(212);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(205)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(205),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => array_obj_ref_672_index_sum_1_req_0); -- 
    -- CP-element group 206 transition  output  bypass 
    -- predecessors 37 
    -- successors 207 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_670_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_670_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_670_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_computed_0
      -- 
    cp_elements(206) <= cp_elements(37);
    index_resize_req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => array_obj_ref_672_index_0_resize_req_0); -- 
    -- CP-element group 207 transition  input  output  no-bypass 
    -- predecessors 206 
    -- successors 208 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resized_0
      -- 
    index_resize_ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_0_resize_ack_0, ack => cp_elements(207)); -- 
    scale_rr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => array_obj_ref_672_index_0_scale_req_0); -- 
    -- CP-element group 208 transition  input  output  no-bypass 
    -- predecessors 207 
    -- successors 209 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_0/scale_ra
      -- 
    scale_ra_2010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_0_scale_ack_0, ack => cp_elements(208)); -- 
    scale_cr_2011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => array_obj_ref_672_index_0_scale_req_1); -- 
    -- CP-element group 209 transition  input  no-bypass 
    -- predecessors 208 
    -- successors 205 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_0/$exit
      -- 
    scale_ca_2012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_0_scale_ack_1, ack => cp_elements(209)); -- 
    -- CP-element group 210 transition  output  bypass 
    -- predecessors 63 
    -- successors 211 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_671_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_671_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_671_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_computed_1
      -- 
    cp_elements(210) <= cp_elements(63);
    index_resize_req_2021_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => array_obj_ref_672_index_1_resize_req_0); -- 
    -- CP-element group 211 transition  input  output  no-bypass 
    -- predecessors 210 
    -- successors 212 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_resized_1
      -- 
    index_resize_ack_2022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_1_resize_ack_0, ack => cp_elements(211)); -- 
    scale_rename_req_2026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => array_obj_ref_672_index_1_rename_req_0); -- 
    -- CP-element group 212 transition  input  no-bypass 
    -- predecessors 211 
    -- successors 205 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_index_scale_1/$exit
      -- 
    scale_rename_ack_2027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_1_rename_ack_0, ack => cp_elements(212)); -- 
    -- CP-element group 213 transition  input  output  no-bypass 
    -- predecessors 205 
    -- successors 214 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_2032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_sum_1_ack_0, ack => cp_elements(213)); -- 
    partial_sum_1_cr_2033_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => array_obj_ref_672_index_sum_1_req_1); -- 
    -- CP-element group 214 transition  input  output  no-bypass 
    -- predecessors 213 
    -- successors 215 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_2034_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_index_sum_1_ack_1, ack => cp_elements(214)); -- 
    final_index_req_2035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(214), ack => array_obj_ref_672_offset_inst_req_0); -- 
    -- CP-element group 215 transition  input  output  no-bypass 
    -- predecessors 214 
    -- successors 216 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_offset_calculated
      -- 
    final_index_ack_2036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_offset_inst_ack_0, ack => cp_elements(215)); -- 
    sum_rename_req_2040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(215), ack => array_obj_ref_672_root_address_inst_req_0); -- 
    -- CP-element group 216 transition  input  no-bypass 
    -- predecessors 215 
    -- successors 203 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_672_root_address_calculated
      -- 
    sum_rename_ack_2041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_672_root_address_inst_ack_0, ack => cp_elements(216)); -- 
    -- CP-element group 217 transition  output  bypass 
    -- predecessors 203 
    -- successors 218 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_673_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_673_complete/$entry
      -- 
    cp_elements(217) <= cp_elements(203);
    final_reg_req_2045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => addr_of_673_final_reg_req_0); -- 
    -- CP-element group 218 transition  input  no-bypass 
    -- predecessors 217 
    -- successors 204 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_673_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_673_complete/$exit
      -- 
    final_reg_ack_2046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_673_final_reg_ack_0, ack => cp_elements(218)); -- 
    -- CP-element group 219 transition  bypass 
    -- predecessors 37 
    -- successors 220 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_679_trigger_
      -- 
    cp_elements(219) <= cp_elements(37);
    -- CP-element group 220 join  fork  transition  bypass 
    -- predecessors 219 233 
    -- successors 221 234 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_679_active_
      -- 
    cpelement_group_220 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(219);
      predecessors(1) <= cp_elements(233);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(220)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(220),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 221 join  transition  no-bypass 
    -- predecessors 220 235 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_679_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_680_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_680_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_680_trigger_
      -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(220);
      predecessors(1) <= cp_elements(235);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(221)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 222 join  transition  output  bypass 
    -- predecessors 226 229 
    -- successors 230 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_indices_scaled
      -- 
    cpelement_group_222 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(226);
      predecessors(1) <= cp_elements(229);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(222)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(222),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => array_obj_ref_678_index_sum_1_req_0); -- 
    -- CP-element group 223 transition  output  bypass 
    -- predecessors 37 
    -- successors 224 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_676_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_676_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_676_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_computed_0
      -- 
    cp_elements(223) <= cp_elements(37);
    index_resize_req_2064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => array_obj_ref_678_index_0_resize_req_0); -- 
    -- CP-element group 224 transition  input  output  no-bypass 
    -- predecessors 223 
    -- successors 225 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resized_0
      -- 
    index_resize_ack_2065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_0_resize_ack_0, ack => cp_elements(224)); -- 
    scale_rr_2069_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => array_obj_ref_678_index_0_scale_req_0); -- 
    -- CP-element group 225 transition  input  output  no-bypass 
    -- predecessors 224 
    -- successors 226 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_0/scale_ra
      -- 
    scale_ra_2070_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_0_scale_ack_0, ack => cp_elements(225)); -- 
    scale_cr_2071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => array_obj_ref_678_index_0_scale_req_1); -- 
    -- CP-element group 226 transition  input  no-bypass 
    -- predecessors 225 
    -- successors 222 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_0/$exit
      -- 
    scale_ca_2072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_0_scale_ack_1, ack => cp_elements(226)); -- 
    -- CP-element group 227 transition  output  bypass 
    -- predecessors 87 
    -- successors 228 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_677_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_677_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_677_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_computed_1
      -- 
    cp_elements(227) <= cp_elements(87);
    index_resize_req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => array_obj_ref_678_index_1_resize_req_0); -- 
    -- CP-element group 228 transition  input  output  no-bypass 
    -- predecessors 227 
    -- successors 229 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_resized_1
      -- 
    index_resize_ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_1_resize_ack_0, ack => cp_elements(228)); -- 
    scale_rename_req_2086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => array_obj_ref_678_index_1_rename_req_0); -- 
    -- CP-element group 229 transition  input  no-bypass 
    -- predecessors 228 
    -- successors 222 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_index_scale_1/$exit
      -- 
    scale_rename_ack_2087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_1_rename_ack_0, ack => cp_elements(229)); -- 
    -- CP-element group 230 transition  input  output  no-bypass 
    -- predecessors 222 
    -- successors 231 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_2092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_sum_1_ack_0, ack => cp_elements(230)); -- 
    partial_sum_1_cr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => array_obj_ref_678_index_sum_1_req_1); -- 
    -- CP-element group 231 transition  input  output  no-bypass 
    -- predecessors 230 
    -- successors 232 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_2094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_index_sum_1_ack_1, ack => cp_elements(231)); -- 
    final_index_req_2095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => array_obj_ref_678_offset_inst_req_0); -- 
    -- CP-element group 232 transition  input  output  no-bypass 
    -- predecessors 231 
    -- successors 233 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_offset_calculated
      -- 
    final_index_ack_2096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_offset_inst_ack_0, ack => cp_elements(232)); -- 
    sum_rename_req_2100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(232), ack => array_obj_ref_678_root_address_inst_req_0); -- 
    -- CP-element group 233 transition  input  no-bypass 
    -- predecessors 232 
    -- successors 220 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_678_root_address_calculated
      -- 
    sum_rename_ack_2101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_678_root_address_inst_ack_0, ack => cp_elements(233)); -- 
    -- CP-element group 234 transition  output  bypass 
    -- predecessors 220 
    -- successors 235 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_679_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_679_complete/$entry
      -- 
    cp_elements(234) <= cp_elements(220);
    final_reg_req_2105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => addr_of_679_final_reg_req_0); -- 
    -- CP-element group 235 transition  input  no-bypass 
    -- predecessors 234 
    -- successors 221 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_679_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_679_complete/$exit
      -- 
    final_reg_ack_2106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_679_final_reg_ack_0, ack => cp_elements(235)); -- 
    -- CP-element group 236 transition  bypass 
    -- predecessors 37 
    -- successors 237 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_685_trigger_
      -- 
    cp_elements(236) <= cp_elements(37);
    -- CP-element group 237 join  fork  transition  bypass 
    -- predecessors 236 250 
    -- successors 238 251 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_685_active_
      -- 
    cpelement_group_237 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(236);
      predecessors(1) <= cp_elements(250);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(237)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(237),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 238 join  transition  no-bypass 
    -- predecessors 237 252 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_685_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_686_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_686_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_686_trigger_
      -- 
    cpelement_group_238 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(237);
      predecessors(1) <= cp_elements(252);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(238)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(238),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 239 join  transition  output  bypass 
    -- predecessors 243 246 
    -- successors 247 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_indices_scaled
      -- 
    cpelement_group_239 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(243);
      predecessors(1) <= cp_elements(246);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(239)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(239),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2151_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => array_obj_ref_684_index_sum_1_req_0); -- 
    -- CP-element group 240 transition  output  bypass 
    -- predecessors 37 
    -- successors 241 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_682_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_682_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_682_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_computed_0
      -- 
    cp_elements(240) <= cp_elements(37);
    index_resize_req_2124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => array_obj_ref_684_index_0_resize_req_0); -- 
    -- CP-element group 241 transition  input  output  no-bypass 
    -- predecessors 240 
    -- successors 242 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resized_0
      -- 
    index_resize_ack_2125_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_index_0_resize_ack_0, ack => cp_elements(241)); -- 
    scale_rr_2129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => array_obj_ref_684_index_0_scale_req_0); -- 
    -- CP-element group 242 transition  input  output  no-bypass 
    -- predecessors 241 
    -- successors 243 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_0/scale_ra
      -- 
    scale_ra_2130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_index_0_scale_ack_0, ack => cp_elements(242)); -- 
    scale_cr_2131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => array_obj_ref_684_index_0_scale_req_1); -- 
    -- CP-element group 243 transition  input  no-bypass 
    -- predecessors 242 
    -- successors 239 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_0/$exit
      -- 
    scale_ca_2132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_index_0_scale_ack_1, ack => cp_elements(243)); -- 
    -- CP-element group 244 transition  output  bypass 
    -- predecessors 162 
    -- successors 245 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_683_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_683_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_683_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_computed_1
      -- 
    cp_elements(244) <= cp_elements(162);
    index_resize_req_2141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => array_obj_ref_684_index_1_resize_req_0); -- 
    -- CP-element group 245 transition  input  output  no-bypass 
    -- predecessors 244 
    -- successors 246 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_resized_1
      -- 
    index_resize_ack_2142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_index_1_resize_ack_0, ack => cp_elements(245)); -- 
    scale_rename_req_2146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(245), ack => array_obj_ref_684_index_1_rename_req_0); -- 
    -- CP-element group 246 transition  input  no-bypass 
    -- predecessors 245 
    -- successors 239 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_index_scale_1/$exit
      -- 
    scale_rename_ack_2147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_index_1_rename_ack_0, ack => cp_elements(246)); -- 
    -- CP-element group 247 transition  input  output  no-bypass 
    -- predecessors 239 
    -- successors 248 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_2152_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_index_sum_1_ack_0, ack => cp_elements(247)); -- 
    partial_sum_1_cr_2153_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(247), ack => array_obj_ref_684_index_sum_1_req_1); -- 
    -- CP-element group 248 transition  input  output  no-bypass 
    -- predecessors 247 
    -- successors 249 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_2154_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_index_sum_1_ack_1, ack => cp_elements(248)); -- 
    final_index_req_2155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => array_obj_ref_684_offset_inst_req_0); -- 
    -- CP-element group 249 transition  input  output  no-bypass 
    -- predecessors 248 
    -- successors 250 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_offset_calculated
      -- 
    final_index_ack_2156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_offset_inst_ack_0, ack => cp_elements(249)); -- 
    sum_rename_req_2160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => array_obj_ref_684_root_address_inst_req_0); -- 
    -- CP-element group 250 transition  input  no-bypass 
    -- predecessors 249 
    -- successors 237 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_684_root_address_calculated
      -- 
    sum_rename_ack_2161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_684_root_address_inst_ack_0, ack => cp_elements(250)); -- 
    -- CP-element group 251 transition  output  bypass 
    -- predecessors 237 
    -- successors 252 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_685_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_685_complete/$entry
      -- 
    cp_elements(251) <= cp_elements(237);
    final_reg_req_2165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => addr_of_685_final_reg_req_0); -- 
    -- CP-element group 252 transition  input  no-bypass 
    -- predecessors 251 
    -- successors 238 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_685_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_685_complete/$exit
      -- 
    final_reg_ack_2166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_685_final_reg_ack_0, ack => cp_elements(252)); -- 
    -- CP-element group 253 transition  bypass 
    -- predecessors 37 
    -- successors 254 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_691_trigger_
      -- 
    cp_elements(253) <= cp_elements(37);
    -- CP-element group 254 join  fork  transition  bypass 
    -- predecessors 253 267 
    -- successors 255 268 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_691_active_
      -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(253);
      predecessors(1) <= cp_elements(267);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(254)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 255 join  transition  no-bypass 
    -- predecessors 254 269 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_691_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_692_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_692_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_692_trigger_
      -- 
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(254);
      predecessors(1) <= cp_elements(269);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(255)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 256 join  transition  output  bypass 
    -- predecessors 260 263 
    -- successors 264 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/$entry
      -- 
    cpelement_group_256 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(260);
      predecessors(1) <= cp_elements(263);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(256)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(256),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => array_obj_ref_690_index_sum_1_req_0); -- 
    -- CP-element group 257 transition  output  bypass 
    -- predecessors 37 
    -- successors 258 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_688_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_688_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_688_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_0/index_resize_req
      -- 
    cp_elements(257) <= cp_elements(37);
    index_resize_req_2184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => array_obj_ref_690_index_0_resize_req_0); -- 
    -- CP-element group 258 transition  input  output  no-bypass 
    -- predecessors 257 
    -- successors 259 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_0/scale_rr
      -- 
    index_resize_ack_2185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_index_0_resize_ack_0, ack => cp_elements(258)); -- 
    scale_rr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => array_obj_ref_690_index_0_scale_req_0); -- 
    -- CP-element group 259 transition  input  output  no-bypass 
    -- predecessors 258 
    -- successors 260 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_0/scale_cr
      -- 
    scale_ra_2190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_index_0_scale_ack_0, ack => cp_elements(259)); -- 
    scale_cr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => array_obj_ref_690_index_0_scale_req_1); -- 
    -- CP-element group 260 transition  input  no-bypass 
    -- predecessors 259 
    -- successors 256 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_0/scale_ca
      -- 
    scale_ca_2192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_index_0_scale_ack_1, ack => cp_elements(260)); -- 
    -- CP-element group 261 transition  output  bypass 
    -- predecessors 39 
    -- successors 262 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_689_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_689_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_689_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_1/index_resize_req
      -- 
    cp_elements(261) <= cp_elements(39);
    index_resize_req_2201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => array_obj_ref_690_index_1_resize_req_0); -- 
    -- CP-element group 262 transition  input  output  no-bypass 
    -- predecessors 261 
    -- successors 263 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_1/$entry
      -- 
    index_resize_ack_2202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_index_1_resize_ack_0, ack => cp_elements(262)); -- 
    scale_rename_req_2206_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(262), ack => array_obj_ref_690_index_1_rename_req_0); -- 
    -- CP-element group 263 transition  input  no-bypass 
    -- predecessors 262 
    -- successors 256 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_index_scale_1/$exit
      -- 
    scale_rename_ack_2207_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_index_1_rename_ack_0, ack => cp_elements(263)); -- 
    -- CP-element group 264 transition  input  output  no-bypass 
    -- predecessors 256 
    -- successors 265 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_2212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_index_sum_1_ack_0, ack => cp_elements(264)); -- 
    partial_sum_1_cr_2213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => array_obj_ref_690_index_sum_1_req_1); -- 
    -- CP-element group 265 transition  input  output  no-bypass 
    -- predecessors 264 
    -- successors 266 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_2214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_index_sum_1_ack_1, ack => cp_elements(265)); -- 
    final_index_req_2215_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => array_obj_ref_690_offset_inst_req_0); -- 
    -- CP-element group 266 transition  input  output  no-bypass 
    -- predecessors 265 
    -- successors 267 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_add_indices/$exit
      -- 
    final_index_ack_2216_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_offset_inst_ack_0, ack => cp_elements(266)); -- 
    sum_rename_req_2220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => array_obj_ref_690_root_address_inst_req_0); -- 
    -- CP-element group 267 transition  input  no-bypass 
    -- predecessors 266 
    -- successors 254 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_690_base_plus_offset/$exit
      -- 
    sum_rename_ack_2221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_690_root_address_inst_ack_0, ack => cp_elements(267)); -- 
    -- CP-element group 268 transition  output  bypass 
    -- predecessors 254 
    -- successors 269 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_691_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_691_complete/final_reg_req
      -- 
    cp_elements(268) <= cp_elements(254);
    final_reg_req_2225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => addr_of_691_final_reg_req_0); -- 
    -- CP-element group 269 transition  input  no-bypass 
    -- predecessors 268 
    -- successors 255 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_691_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_691_complete/$exit
      -- 
    final_reg_ack_2226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_691_final_reg_ack_0, ack => cp_elements(269)); -- 
    -- CP-element group 270 transition  bypass 
    -- predecessors 37 
    -- successors 271 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_697_trigger_
      -- 
    cp_elements(270) <= cp_elements(37);
    -- CP-element group 271 join  fork  transition  bypass 
    -- predecessors 270 284 
    -- successors 272 285 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_697_active_
      -- 
    cpelement_group_271 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(270);
      predecessors(1) <= cp_elements(284);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(271)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(271),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 272 join  transition  no-bypass 
    -- predecessors 271 286 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_698_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_697_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_698_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_698_completed_
      -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(271);
      predecessors(1) <= cp_elements(286);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(272)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 273 join  transition  output  bypass 
    -- predecessors 277 280 
    -- successors 281 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/$entry
      -- 
    cpelement_group_273 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(277);
      predecessors(1) <= cp_elements(280);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(273)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(273),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => array_obj_ref_696_index_sum_1_req_0); -- 
    -- CP-element group 274 transition  output  bypass 
    -- predecessors 37 
    -- successors 275 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_694_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_694_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_694_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_0/$entry
      -- 
    cp_elements(274) <= cp_elements(37);
    index_resize_req_2244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => array_obj_ref_696_index_0_resize_req_0); -- 
    -- CP-element group 275 transition  input  output  no-bypass 
    -- predecessors 274 
    -- successors 276 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_0/$exit
      -- 
    index_resize_ack_2245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_index_0_resize_ack_0, ack => cp_elements(275)); -- 
    scale_rr_2249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => array_obj_ref_696_index_0_scale_req_0); -- 
    -- CP-element group 276 transition  input  output  no-bypass 
    -- predecessors 275 
    -- successors 277 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_0/scale_cr
      -- 
    scale_ra_2250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_index_0_scale_ack_0, ack => cp_elements(276)); -- 
    scale_cr_2251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(276), ack => array_obj_ref_696_index_0_scale_req_1); -- 
    -- CP-element group 277 transition  input  no-bypass 
    -- predecessors 276 
    -- successors 273 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_0/$exit
      -- 
    scale_ca_2252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_index_0_scale_ack_1, ack => cp_elements(277)); -- 
    -- CP-element group 278 transition  output  bypass 
    -- predecessors 63 
    -- successors 279 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_695_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_695_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_695_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_1/index_resize_req
      -- 
    cp_elements(278) <= cp_elements(63);
    index_resize_req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(278), ack => array_obj_ref_696_index_1_resize_req_0); -- 
    -- CP-element group 279 transition  input  output  no-bypass 
    -- predecessors 278 
    -- successors 280 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_index_1_resize_ack_0, ack => cp_elements(279)); -- 
    scale_rename_req_2266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => array_obj_ref_696_index_1_rename_req_0); -- 
    -- CP-element group 280 transition  input  no-bypass 
    -- predecessors 279 
    -- successors 273 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_index_scale_1/$exit
      -- 
    scale_rename_ack_2267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_index_1_rename_ack_0, ack => cp_elements(280)); -- 
    -- CP-element group 281 transition  input  output  no-bypass 
    -- predecessors 273 
    -- successors 282 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_2272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_index_sum_1_ack_0, ack => cp_elements(281)); -- 
    partial_sum_1_cr_2273_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(281), ack => array_obj_ref_696_index_sum_1_req_1); -- 
    -- CP-element group 282 transition  input  output  no-bypass 
    -- predecessors 281 
    -- successors 283 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2274_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_index_sum_1_ack_1, ack => cp_elements(282)); -- 
    final_index_req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => array_obj_ref_696_offset_inst_req_0); -- 
    -- CP-element group 283 transition  input  output  no-bypass 
    -- predecessors 282 
    -- successors 284 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_add_indices/$exit
      -- 
    final_index_ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_offset_inst_ack_0, ack => cp_elements(283)); -- 
    sum_rename_req_2280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(283), ack => array_obj_ref_696_root_address_inst_req_0); -- 
    -- CP-element group 284 transition  input  no-bypass 
    -- predecessors 283 
    -- successors 271 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_696_root_address_calculated
      -- 
    sum_rename_ack_2281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_696_root_address_inst_ack_0, ack => cp_elements(284)); -- 
    -- CP-element group 285 transition  output  bypass 
    -- predecessors 271 
    -- successors 286 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_697_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_697_complete/final_reg_req
      -- 
    cp_elements(285) <= cp_elements(271);
    final_reg_req_2285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(285), ack => addr_of_697_final_reg_req_0); -- 
    -- CP-element group 286 transition  input  no-bypass 
    -- predecessors 285 
    -- successors 272 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_697_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_697_complete/final_reg_ack
      -- 
    final_reg_ack_2286_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_697_final_reg_ack_0, ack => cp_elements(286)); -- 
    -- CP-element group 287 transition  bypass 
    -- predecessors 37 
    -- successors 288 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_703_trigger_
      -- 
    cp_elements(287) <= cp_elements(37);
    -- CP-element group 288 join  fork  transition  bypass 
    -- predecessors 287 301 
    -- successors 289 302 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_703_active_
      -- 
    cpelement_group_288 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(287);
      predecessors(1) <= cp_elements(301);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(288)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(288),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 289 join  transition  no-bypass 
    -- predecessors 288 303 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_704_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_704_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_704_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_703_completed_
      -- 
    cpelement_group_289 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(288);
      predecessors(1) <= cp_elements(303);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(289)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(289),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 290 join  transition  output  bypass 
    -- predecessors 294 297 
    -- successors 298 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_indices_scaled
      -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(294);
      predecessors(1) <= cp_elements(297);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(290)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => array_obj_ref_702_index_sum_1_req_0); -- 
    -- CP-element group 291 transition  output  bypass 
    -- predecessors 37 
    -- successors 292 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_700_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_700_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_700_active_
      -- 
    cp_elements(291) <= cp_elements(37);
    index_resize_req_2304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(291), ack => array_obj_ref_702_index_0_resize_req_0); -- 
    -- CP-element group 292 transition  input  output  no-bypass 
    -- predecessors 291 
    -- successors 293 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_index_0_resize_ack_0, ack => cp_elements(292)); -- 
    scale_rr_2309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => array_obj_ref_702_index_0_scale_req_0); -- 
    -- CP-element group 293 transition  input  output  no-bypass 
    -- predecessors 292 
    -- successors 294 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_0/scale_cr
      -- 
    scale_ra_2310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_index_0_scale_ack_0, ack => cp_elements(293)); -- 
    scale_cr_2311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(293), ack => array_obj_ref_702_index_0_scale_req_1); -- 
    -- CP-element group 294 transition  input  no-bypass 
    -- predecessors 293 
    -- successors 290 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_0/scale_ca
      -- 
    scale_ca_2312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_index_0_scale_ack_1, ack => cp_elements(294)); -- 
    -- CP-element group 295 transition  output  bypass 
    -- predecessors 87 
    -- successors 296 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_701_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_701_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_701_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_1/index_resize_req
      -- 
    cp_elements(295) <= cp_elements(87);
    index_resize_req_2321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(295), ack => array_obj_ref_702_index_1_resize_req_0); -- 
    -- CP-element group 296 transition  input  output  no-bypass 
    -- predecessors 295 
    -- successors 297 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_index_1_resize_ack_0, ack => cp_elements(296)); -- 
    scale_rename_req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(296), ack => array_obj_ref_702_index_1_rename_req_0); -- 
    -- CP-element group 297 transition  input  no-bypass 
    -- predecessors 296 
    -- successors 290 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_index_1_rename_ack_0, ack => cp_elements(297)); -- 
    -- CP-element group 298 transition  input  output  no-bypass 
    -- predecessors 290 
    -- successors 299 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_2332_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_index_sum_1_ack_0, ack => cp_elements(298)); -- 
    partial_sum_1_cr_2333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => array_obj_ref_702_index_sum_1_req_1); -- 
    -- CP-element group 299 transition  input  output  no-bypass 
    -- predecessors 298 
    -- successors 300 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_index_sum_1_ack_1, ack => cp_elements(299)); -- 
    final_index_req_2335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(299), ack => array_obj_ref_702_offset_inst_req_0); -- 
    -- CP-element group 300 transition  input  output  no-bypass 
    -- predecessors 299 
    -- successors 301 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_offset_calculated
      -- 
    final_index_ack_2336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_offset_inst_ack_0, ack => cp_elements(300)); -- 
    sum_rename_req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => array_obj_ref_702_root_address_inst_req_0); -- 
    -- CP-element group 301 transition  input  no-bypass 
    -- predecessors 300 
    -- successors 288 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_702_root_address_calculated
      -- 
    sum_rename_ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_702_root_address_inst_ack_0, ack => cp_elements(301)); -- 
    -- CP-element group 302 transition  output  bypass 
    -- predecessors 288 
    -- successors 303 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_703_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_703_complete/$entry
      -- 
    cp_elements(302) <= cp_elements(288);
    final_reg_req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(302), ack => addr_of_703_final_reg_req_0); -- 
    -- CP-element group 303 transition  input  no-bypass 
    -- predecessors 302 
    -- successors 289 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_703_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_703_complete/$exit
      -- 
    final_reg_ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_703_final_reg_ack_0, ack => cp_elements(303)); -- 
    -- CP-element group 304 transition  bypass 
    -- predecessors 37 
    -- successors 305 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_709_trigger_
      -- 
    cp_elements(304) <= cp_elements(37);
    -- CP-element group 305 join  fork  transition  bypass 
    -- predecessors 304 318 
    -- successors 306 319 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_709_active_
      -- 
    cpelement_group_305 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(304);
      predecessors(1) <= cp_elements(318);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(305)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(305),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 306 join  transition  no-bypass 
    -- predecessors 305 320 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_710_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_710_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_710_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_709_completed_
      -- 
    cpelement_group_306 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(305);
      predecessors(1) <= cp_elements(320);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(306)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(306),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 307 join  transition  output  bypass 
    -- predecessors 311 314 
    -- successors 315 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_indices_scaled
      -- 
    cpelement_group_307 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(311);
      predecessors(1) <= cp_elements(314);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(307)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(307),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(307), ack => array_obj_ref_708_index_sum_1_req_0); -- 
    -- CP-element group 308 transition  output  bypass 
    -- predecessors 37 
    -- successors 309 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_706_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_706_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_706_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_computed_0
      -- 
    cp_elements(308) <= cp_elements(37);
    index_resize_req_2364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => array_obj_ref_708_index_0_resize_req_0); -- 
    -- CP-element group 309 transition  input  output  no-bypass 
    -- predecessors 308 
    -- successors 310 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resized_0
      -- 
    index_resize_ack_2365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_0_resize_ack_0, ack => cp_elements(309)); -- 
    scale_rr_2369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(309), ack => array_obj_ref_708_index_0_scale_req_0); -- 
    -- CP-element group 310 transition  input  output  no-bypass 
    -- predecessors 309 
    -- successors 311 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_0/scale_cr
      -- 
    scale_ra_2370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_0_scale_ack_0, ack => cp_elements(310)); -- 
    scale_cr_2371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(310), ack => array_obj_ref_708_index_0_scale_req_1); -- 
    -- CP-element group 311 transition  input  no-bypass 
    -- predecessors 310 
    -- successors 307 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_0/$exit
      -- 
    scale_ca_2372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_0_scale_ack_1, ack => cp_elements(311)); -- 
    -- CP-element group 312 transition  output  bypass 
    -- predecessors 162 
    -- successors 313 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_707_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_707_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_707_completed_
      -- 
    cp_elements(312) <= cp_elements(162);
    index_resize_req_2381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(312), ack => array_obj_ref_708_index_1_resize_req_0); -- 
    -- CP-element group 313 transition  input  output  no-bypass 
    -- predecessors 312 
    -- successors 314 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_resize_1/index_resize_ack
      -- 
    index_resize_ack_2382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_1_resize_ack_0, ack => cp_elements(313)); -- 
    scale_rename_req_2386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(313), ack => array_obj_ref_708_index_1_rename_req_0); -- 
    -- CP-element group 314 transition  input  no-bypass 
    -- predecessors 313 
    -- successors 307 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_1_rename_ack_0, ack => cp_elements(314)); -- 
    -- CP-element group 315 transition  input  output  no-bypass 
    -- predecessors 307 
    -- successors 316 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_2392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_sum_1_ack_0, ack => cp_elements(315)); -- 
    partial_sum_1_cr_2393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => array_obj_ref_708_index_sum_1_req_1); -- 
    -- CP-element group 316 transition  input  output  no-bypass 
    -- predecessors 315 
    -- successors 317 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_2394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_index_sum_1_ack_1, ack => cp_elements(316)); -- 
    final_index_req_2395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(316), ack => array_obj_ref_708_offset_inst_req_0); -- 
    -- CP-element group 317 transition  input  output  no-bypass 
    -- predecessors 316 
    -- successors 318 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_add_indices/$exit
      -- 
    final_index_ack_2396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_offset_inst_ack_0, ack => cp_elements(317)); -- 
    sum_rename_req_2400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(317), ack => array_obj_ref_708_root_address_inst_req_0); -- 
    -- CP-element group 318 transition  input  no-bypass 
    -- predecessors 317 
    -- successors 305 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_708_root_address_calculated
      -- 
    sum_rename_ack_2401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_708_root_address_inst_ack_0, ack => cp_elements(318)); -- 
    -- CP-element group 319 transition  output  bypass 
    -- predecessors 305 
    -- successors 320 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_709_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_709_complete/$entry
      -- 
    cp_elements(319) <= cp_elements(305);
    final_reg_req_2405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => addr_of_709_final_reg_req_0); -- 
    -- CP-element group 320 transition  input  no-bypass 
    -- predecessors 319 
    -- successors 306 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_709_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_709_complete/$exit
      -- 
    final_reg_ack_2406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_709_final_reg_ack_0, ack => cp_elements(320)); -- 
    -- CP-element group 321 transition  bypass 
    -- predecessors 37 
    -- successors 322 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_715_trigger_
      -- 
    cp_elements(321) <= cp_elements(37);
    -- CP-element group 322 join  fork  transition  bypass 
    -- predecessors 321 335 
    -- successors 323 336 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_715_active_
      -- 
    cpelement_group_322 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(321);
      predecessors(1) <= cp_elements(335);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(322)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(322),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 323 join  transition  no-bypass 
    -- predecessors 322 337 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_716_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_716_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_716_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_715_completed_
      -- 
    cpelement_group_323 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(322);
      predecessors(1) <= cp_elements(337);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(323)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(323),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 324 join  transition  output  bypass 
    -- predecessors 328 331 
    -- successors 332 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_indices_scaled
      -- 
    cpelement_group_324 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(328);
      predecessors(1) <= cp_elements(331);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(324)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(324),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(324), ack => array_obj_ref_714_index_sum_1_req_0); -- 
    -- CP-element group 325 transition  output  bypass 
    -- predecessors 37 
    -- successors 326 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_712_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_712_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_712_completed_
      -- 
    cp_elements(325) <= cp_elements(37);
    index_resize_req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => array_obj_ref_714_index_0_resize_req_0); -- 
    -- CP-element group 326 transition  input  output  no-bypass 
    -- predecessors 325 
    -- successors 327 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_0/$entry
      -- 
    index_resize_ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_index_0_resize_ack_0, ack => cp_elements(326)); -- 
    scale_rr_2429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(326), ack => array_obj_ref_714_index_0_scale_req_0); -- 
    -- CP-element group 327 transition  input  output  no-bypass 
    -- predecessors 326 
    -- successors 328 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_0/scale_ra
      -- 
    scale_ra_2430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_index_0_scale_ack_0, ack => cp_elements(327)); -- 
    scale_cr_2431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(327), ack => array_obj_ref_714_index_0_scale_req_1); -- 
    -- CP-element group 328 transition  input  no-bypass 
    -- predecessors 327 
    -- successors 324 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_0/$exit
      -- 
    scale_ca_2432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_index_0_scale_ack_1, ack => cp_elements(328)); -- 
    -- CP-element group 329 transition  output  bypass 
    -- predecessors 162 
    -- successors 330 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_713_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_713_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_713_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_1/$entry
      -- 
    cp_elements(329) <= cp_elements(162);
    index_resize_req_2441_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(329), ack => array_obj_ref_714_index_1_resize_req_0); -- 
    -- CP-element group 330 transition  input  output  no-bypass 
    -- predecessors 329 
    -- successors 331 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_resize_1/$exit
      -- 
    index_resize_ack_2442_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_index_1_resize_ack_0, ack => cp_elements(330)); -- 
    scale_rename_req_2446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(330), ack => array_obj_ref_714_index_1_rename_req_0); -- 
    -- CP-element group 331 transition  input  no-bypass 
    -- predecessors 330 
    -- successors 324 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_index_scale_1/$exit
      -- 
    scale_rename_ack_2447_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_index_1_rename_ack_0, ack => cp_elements(331)); -- 
    -- CP-element group 332 transition  input  output  no-bypass 
    -- predecessors 324 
    -- successors 333 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_2452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_index_sum_1_ack_0, ack => cp_elements(332)); -- 
    partial_sum_1_cr_2453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(332), ack => array_obj_ref_714_index_sum_1_req_1); -- 
    -- CP-element group 333 transition  input  output  no-bypass 
    -- predecessors 332 
    -- successors 334 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_index_sum_1_ack_1, ack => cp_elements(333)); -- 
    final_index_req_2455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => array_obj_ref_714_offset_inst_req_0); -- 
    -- CP-element group 334 transition  input  output  no-bypass 
    -- predecessors 333 
    -- successors 335 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_base_plus_offset/$entry
      -- 
    final_index_ack_2456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_offset_inst_ack_0, ack => cp_elements(334)); -- 
    sum_rename_req_2460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(334), ack => array_obj_ref_714_root_address_inst_req_0); -- 
    -- CP-element group 335 transition  input  no-bypass 
    -- predecessors 334 
    -- successors 322 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/array_obj_ref_714_root_address_calculated
      -- 
    sum_rename_ack_2461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_714_root_address_inst_ack_0, ack => cp_elements(335)); -- 
    -- CP-element group 336 transition  output  bypass 
    -- predecessors 322 
    -- successors 337 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_715_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_715_complete/$entry
      -- 
    cp_elements(336) <= cp_elements(322);
    final_reg_req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => addr_of_715_final_reg_req_0); -- 
    -- CP-element group 337 transition  input  no-bypass 
    -- predecessors 336 
    -- successors 323 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_715_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/addr_of_715_complete/$exit
      -- 
    final_reg_ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_715_final_reg_ack_0, ack => cp_elements(337)); -- 
    -- CP-element group 338 join  fork  transition  bypass 
    -- predecessors 340 342 
    -- successors 339 343 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_active_
      -- 
    cpelement_group_338 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(340);
      predecessors(1) <= cp_elements(342);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(338)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(338),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 339 join  fork  transition  no-bypass 
    -- predecessors 338 344 
    -- successors 347 354 361 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_722_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_722_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_722_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_completed_
      -- 
    cpelement_group_339 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(338);
      predecessors(1) <= cp_elements(344);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(339)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(339),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 340 fork  transition  bypass 
    -- predecessors 37 
    -- successors 338 341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_718_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_718_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_718_completed_
      -- 
    cp_elements(340) <= cp_elements(37);
    -- CP-element group 341 transition  output  bypass 
    -- predecessors 340 
    -- successors 342 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Sample/rr
      -- 
    cp_elements(341) <= cp_elements(340);
    rr_2479_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => binary_721_inst_req_0); -- 
    -- CP-element group 342 transition  input  no-bypass 
    -- predecessors 341 
    -- successors 338 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Sample/$exit
      -- 
    ra_2480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_721_inst_ack_0, ack => cp_elements(342)); -- 
    -- CP-element group 343 transition  output  bypass 
    -- predecessors 338 
    -- successors 344 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Update/cr
      -- 
    cp_elements(343) <= cp_elements(338);
    cr_2484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(343), ack => binary_721_inst_req_1); -- 
    -- CP-element group 344 transition  input  no-bypass 
    -- predecessors 343 
    -- successors 339 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_721_complete_Update/ca
      -- 
    ca_2485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_721_inst_ack_1, ack => cp_elements(344)); -- 
    -- CP-element group 345 join  fork  transition  no-bypass 
    -- predecessors 347 349 
    -- successors 346 350 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_active_
      -- 
    cpelement_group_345 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(347);
      predecessors(1) <= cp_elements(349);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(345)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(345),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 346 join  transition  no-bypass 
    -- predecessors 345 351 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_728_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_728_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_728_trigger_
      -- 
    cpelement_group_346 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(345);
      predecessors(1) <= cp_elements(351);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(346)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(346),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 347 fork  transition  bypass 
    -- predecessors 339 
    -- successors 345 348 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_724_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_724_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_724_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_trigger_
      -- 
    cp_elements(347) <= cp_elements(339);
    -- CP-element group 348 transition  output  bypass 
    -- predecessors 347 
    -- successors 349 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Sample/$entry
      -- 
    cp_elements(348) <= cp_elements(347);
    rr_2498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => binary_727_inst_req_0); -- 
    -- CP-element group 349 transition  input  no-bypass 
    -- predecessors 348 
    -- successors 345 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Sample/$exit
      -- 
    ra_2499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_727_inst_ack_0, ack => cp_elements(349)); -- 
    -- CP-element group 350 transition  output  bypass 
    -- predecessors 345 
    -- successors 351 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Update/cr
      -- 
    cp_elements(350) <= cp_elements(345);
    cr_2503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => binary_727_inst_req_1); -- 
    -- CP-element group 351 transition  input  no-bypass 
    -- predecessors 350 
    -- successors 346 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_727_complete_Update/ca
      -- 
    ca_2504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_727_inst_ack_1, ack => cp_elements(351)); -- 
    -- CP-element group 352 join  fork  transition  no-bypass 
    -- predecessors 354 356 
    -- successors 353 357 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_active_
      -- 
    cpelement_group_352 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(354);
      predecessors(1) <= cp_elements(356);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(352)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(352),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 353 join  transition  no-bypass 
    -- predecessors 352 358 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_734_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_734_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_734_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_completed_
      -- 
    cpelement_group_353 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(352);
      predecessors(1) <= cp_elements(358);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(353)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(353),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 354 fork  transition  bypass 
    -- predecessors 339 
    -- successors 352 355 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_730_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_730_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_730_completed_
      -- 
    cp_elements(354) <= cp_elements(339);
    -- CP-element group 355 transition  output  bypass 
    -- predecessors 354 
    -- successors 356 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Sample/rr
      -- 
    cp_elements(355) <= cp_elements(354);
    rr_2517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(355), ack => binary_733_inst_req_0); -- 
    -- CP-element group 356 transition  input  no-bypass 
    -- predecessors 355 
    -- successors 352 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Sample/ra
      -- 
    ra_2518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_733_inst_ack_0, ack => cp_elements(356)); -- 
    -- CP-element group 357 transition  output  bypass 
    -- predecessors 352 
    -- successors 358 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Update/cr
      -- 
    cp_elements(357) <= cp_elements(352);
    cr_2522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => binary_733_inst_req_1); -- 
    -- CP-element group 358 transition  input  no-bypass 
    -- predecessors 357 
    -- successors 353 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_733_complete_Update/ca
      -- 
    ca_2523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_733_inst_ack_1, ack => cp_elements(358)); -- 
    -- CP-element group 359 join  fork  transition  no-bypass 
    -- predecessors 361 363 
    -- successors 360 364 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_active_
      -- 
    cpelement_group_359 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(361);
      predecessors(1) <= cp_elements(363);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(359)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(359),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 360 join  transition  no-bypass 
    -- predecessors 359 365 
    -- successors 366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_740_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_740_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/assign_stmt_740_completed_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_completed_
      -- 
    cpelement_group_360 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(359);
      predecessors(1) <= cp_elements(365);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(360)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(360),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 361 fork  transition  bypass 
    -- predecessors 339 
    -- successors 359 362 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_736_trigger_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_736_active_
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/simple_obj_ref_736_completed_
      -- 
    cp_elements(361) <= cp_elements(339);
    -- CP-element group 362 transition  output  bypass 
    -- predecessors 361 
    -- successors 363 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Sample/rr
      -- 
    cp_elements(362) <= cp_elements(361);
    rr_2536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(362), ack => binary_739_inst_req_0); -- 
    -- CP-element group 363 transition  input  no-bypass 
    -- predecessors 362 
    -- successors 359 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Sample/ra
      -- 
    ra_2537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_739_inst_ack_0, ack => cp_elements(363)); -- 
    -- CP-element group 364 transition  output  bypass 
    -- predecessors 359 
    -- successors 365 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Update/cr
      -- 
    cp_elements(364) <= cp_elements(359);
    cr_2541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(364), ack => binary_739_inst_req_1); -- 
    -- CP-element group 365 transition  input  no-bypass 
    -- predecessors 364 
    -- successors 360 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/binary_739_complete_Update/ca
      -- 
    ca_2542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_739_inst_ack_1, ack => cp_elements(365)); -- 
    -- CP-element group 366 join  transition  bypass 
    -- predecessors 47 71 95 112 129 146 170 187 204 221 238 255 272 289 306 323 346 353 360 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740/$exit
      -- 
    cpelement_group_366 : Block -- 
      signal predecessors: BooleanArray(18 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(47);
      predecessors(1) <= cp_elements(71);
      predecessors(2) <= cp_elements(95);
      predecessors(3) <= cp_elements(112);
      predecessors(4) <= cp_elements(129);
      predecessors(5) <= cp_elements(146);
      predecessors(6) <= cp_elements(170);
      predecessors(7) <= cp_elements(187);
      predecessors(8) <= cp_elements(204);
      predecessors(9) <= cp_elements(221);
      predecessors(10) <= cp_elements(238);
      predecessors(11) <= cp_elements(255);
      predecessors(12) <= cp_elements(272);
      predecessors(13) <= cp_elements(289);
      predecessors(14) <= cp_elements(306);
      predecessors(15) <= cp_elements(323);
      predecessors(16) <= cp_elements(346);
      predecessors(17) <= cp_elements(353);
      predecessors(18) <= cp_elements(360);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(366)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(366),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 367 fork  transition  bypass 
    -- predecessors 3 
    -- successors 370 375 379 399 403 423 427 440 444 457 461 474 478 498 502 515 519 532 536 549 553 566 570 583 587 600 604 617 621 634 638 651 655 670 682 690 706 714 730 738 747 755 764 772 781 789 798 806 815 823 832 840 849 857 866 874 883 891 900 908 917 925 934 942 951 959 1108 1213 1318 1423 1528 1593 1658 1723 1828 1893 1958 2023 2128 2193 2258 2323 2330 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/$entry
      -- 
    cp_elements(367) <= cp_elements(3);
    -- CP-element group 368 join  fork  transition  no-bypass 
    -- predecessors 370 372 
    -- successors 369 373 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_active_
      -- 
    cpelement_group_368 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(370);
      predecessors(1) <= cp_elements(372);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(368)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(368),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 369 join  fork  transition  bypass 
    -- predecessors 368 374 
    -- successors 383 394 418 448 493 523 591 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_868_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_868_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_868_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_completed_
      -- 
    cpelement_group_369 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(368);
      predecessors(1) <= cp_elements(374);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(369)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(369),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 370 fork  transition  bypass 
    -- predecessors 367 
    -- successors 368 371 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_864_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_864_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_864_completed_
      -- 
    cp_elements(370) <= cp_elements(367);
    -- CP-element group 371 transition  output  bypass 
    -- predecessors 370 
    -- successors 372 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Sample/rr
      -- 
    cp_elements(371) <= cp_elements(370);
    rr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(371), ack => binary_867_inst_req_0); -- 
    -- CP-element group 372 transition  input  no-bypass 
    -- predecessors 371 
    -- successors 368 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Sample/ra
      -- 
    ra_2559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_867_inst_ack_0, ack => cp_elements(372)); -- 
    -- CP-element group 373 transition  output  bypass 
    -- predecessors 368 
    -- successors 374 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Update/cr
      -- 
    cp_elements(373) <= cp_elements(368);
    cr_2563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(373), ack => binary_867_inst_req_1); -- 
    -- CP-element group 374 transition  input  no-bypass 
    -- predecessors 373 
    -- successors 369 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_867_complete_Update/ca
      -- 
    ca_2564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_867_inst_ack_1, ack => cp_elements(374)); -- 
    -- CP-element group 375 transition  bypass 
    -- predecessors 367 
    -- successors 376 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_873_trigger_
      -- 
    cp_elements(375) <= cp_elements(367);
    -- CP-element group 376 join  fork  transition  no-bypass 
    -- predecessors 375 389 
    -- successors 377 390 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_873_active_
      -- 
    cpelement_group_376 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(375);
      predecessors(1) <= cp_elements(389);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(376)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(376),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 377 join  transition  output  bypass 
    -- predecessors 376 391 
    -- successors 970 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_874_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_874_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_874_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_873_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1104_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1104_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1104_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_addr_resize/base_resize_req
      -- 
    cpelement_group_377 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(376);
      predecessors(1) <= cp_elements(391);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(377)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(377),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(377), ack => ptr_deref_1105_base_resize_req_0); -- 
    -- CP-element group 378 join  transition  output  bypass 
    -- predecessors 382 385 
    -- successors 386 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_378 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(382);
      predecessors(1) <= cp_elements(385);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(378)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(378),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(378), ack => array_obj_ref_872_index_sum_1_req_0); -- 
    -- CP-element group 379 transition  output  bypass 
    -- predecessors 367 
    -- successors 380 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_870_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_870_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_870_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_0/index_resize_req
      -- 
    cp_elements(379) <= cp_elements(367);
    index_resize_req_2582_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(379), ack => array_obj_ref_872_index_0_resize_req_0); -- 
    -- CP-element group 380 transition  input  output  no-bypass 
    -- predecessors 379 
    -- successors 381 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_0/scale_rr
      -- 
    index_resize_ack_2583_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_index_0_resize_ack_0, ack => cp_elements(380)); -- 
    scale_rr_2587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => array_obj_ref_872_index_0_scale_req_0); -- 
    -- CP-element group 381 transition  input  output  no-bypass 
    -- predecessors 380 
    -- successors 382 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_0/scale_cr
      -- 
    scale_ra_2588_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_index_0_scale_ack_0, ack => cp_elements(381)); -- 
    scale_cr_2589_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => array_obj_ref_872_index_0_scale_req_1); -- 
    -- CP-element group 382 transition  input  no-bypass 
    -- predecessors 381 
    -- successors 378 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_0/scale_ca
      -- 
    scale_ca_2590_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_index_0_scale_ack_1, ack => cp_elements(382)); -- 
    -- CP-element group 383 transition  output  bypass 
    -- predecessors 369 
    -- successors 384 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_871_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_871_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_871_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_1/index_resize_req
      -- 
    cp_elements(383) <= cp_elements(369);
    index_resize_req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(383), ack => array_obj_ref_872_index_1_resize_req_0); -- 
    -- CP-element group 384 transition  input  output  no-bypass 
    -- predecessors 383 
    -- successors 385 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_index_1_resize_ack_0, ack => cp_elements(384)); -- 
    scale_rename_req_2604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(384), ack => array_obj_ref_872_index_1_rename_req_0); -- 
    -- CP-element group 385 transition  input  no-bypass 
    -- predecessors 384 
    -- successors 378 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_index_1_rename_ack_0, ack => cp_elements(385)); -- 
    -- CP-element group 386 transition  input  output  no-bypass 
    -- predecessors 378 
    -- successors 387 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_2610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_index_sum_1_ack_0, ack => cp_elements(386)); -- 
    partial_sum_1_cr_2611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(386), ack => array_obj_ref_872_index_sum_1_req_1); -- 
    -- CP-element group 387 transition  input  output  no-bypass 
    -- predecessors 386 
    -- successors 388 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_index_sum_1_ack_1, ack => cp_elements(387)); -- 
    final_index_req_2613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(387), ack => array_obj_ref_872_offset_inst_req_0); -- 
    -- CP-element group 388 transition  input  output  no-bypass 
    -- predecessors 387 
    -- successors 389 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_2614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_offset_inst_ack_0, ack => cp_elements(388)); -- 
    sum_rename_req_2618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(388), ack => array_obj_ref_872_root_address_inst_req_0); -- 
    -- CP-element group 389 transition  input  no-bypass 
    -- predecessors 388 
    -- successors 376 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_872_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_872_root_address_inst_ack_0, ack => cp_elements(389)); -- 
    -- CP-element group 390 transition  output  bypass 
    -- predecessors 376 
    -- successors 391 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_873_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_873_complete/final_reg_req
      -- 
    cp_elements(390) <= cp_elements(376);
    final_reg_req_2623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(390), ack => addr_of_873_final_reg_req_0); -- 
    -- CP-element group 391 transition  input  no-bypass 
    -- predecessors 390 
    -- successors 377 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_873_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_873_complete/final_reg_ack
      -- 
    final_reg_ack_2624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_873_final_reg_ack_0, ack => cp_elements(391)); -- 
    -- CP-element group 392 join  fork  transition  no-bypass 
    -- predecessors 394 396 
    -- successors 393 397 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_active_
      -- 
    cpelement_group_392 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(394);
      predecessors(1) <= cp_elements(396);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(392)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(392),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 393 join  fork  transition  no-bypass 
    -- predecessors 392 398 
    -- successors 407 465 540 608 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_880_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_880_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_880_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_completed_
      -- 
    cpelement_group_393 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(392);
      predecessors(1) <= cp_elements(398);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(393)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(393),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 394 fork  transition  bypass 
    -- predecessors 369 
    -- successors 392 395 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_876_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_876_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_876_completed_
      -- 
    cp_elements(394) <= cp_elements(369);
    -- CP-element group 395 transition  output  bypass 
    -- predecessors 394 
    -- successors 396 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Sample/rr
      -- 
    cp_elements(395) <= cp_elements(394);
    rr_2637_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(395), ack => binary_879_inst_req_0); -- 
    -- CP-element group 396 transition  input  no-bypass 
    -- predecessors 395 
    -- successors 392 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Sample/ra
      -- 
    ra_2638_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_879_inst_ack_0, ack => cp_elements(396)); -- 
    -- CP-element group 397 transition  output  bypass 
    -- predecessors 392 
    -- successors 398 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Update/cr
      -- 
    cp_elements(397) <= cp_elements(392);
    cr_2642_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(397), ack => binary_879_inst_req_1); -- 
    -- CP-element group 398 transition  input  no-bypass 
    -- predecessors 397 
    -- successors 393 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_879_complete_Update/ca
      -- 
    ca_2643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_879_inst_ack_1, ack => cp_elements(398)); -- 
    -- CP-element group 399 transition  bypass 
    -- predecessors 367 
    -- successors 400 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_885_trigger_
      -- 
    cp_elements(399) <= cp_elements(367);
    -- CP-element group 400 join  fork  transition  no-bypass 
    -- predecessors 399 413 
    -- successors 401 414 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_885_active_
      -- 
    cpelement_group_400 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(399);
      predecessors(1) <= cp_elements(413);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(400)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(400),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 401 join  transition  output  bypass 
    -- predecessors 400 415 
    -- successors 1030 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_886_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_886_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_886_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_885_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1128_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1128_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1128_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_addr_resize/base_resize_req
      -- 
    cpelement_group_401 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(400);
      predecessors(1) <= cp_elements(415);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(401)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(401),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4946_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(401), ack => ptr_deref_1129_base_resize_req_0); -- 
    -- CP-element group 402 join  transition  output  bypass 
    -- predecessors 406 409 
    -- successors 410 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_402 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(406);
      predecessors(1) <= cp_elements(409);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(402)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(402),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(402), ack => array_obj_ref_884_index_sum_1_req_0); -- 
    -- CP-element group 403 transition  output  bypass 
    -- predecessors 367 
    -- successors 404 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_882_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_882_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_882_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_0/index_resize_req
      -- 
    cp_elements(403) <= cp_elements(367);
    index_resize_req_2661_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(403), ack => array_obj_ref_884_index_0_resize_req_0); -- 
    -- CP-element group 404 transition  input  output  no-bypass 
    -- predecessors 403 
    -- successors 405 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_0/scale_rr
      -- 
    index_resize_ack_2662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_0_resize_ack_0, ack => cp_elements(404)); -- 
    scale_rr_2666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(404), ack => array_obj_ref_884_index_0_scale_req_0); -- 
    -- CP-element group 405 transition  input  output  no-bypass 
    -- predecessors 404 
    -- successors 406 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_0/scale_cr
      -- 
    scale_ra_2667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_0_scale_ack_0, ack => cp_elements(405)); -- 
    scale_cr_2668_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(405), ack => array_obj_ref_884_index_0_scale_req_1); -- 
    -- CP-element group 406 transition  input  no-bypass 
    -- predecessors 405 
    -- successors 402 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_0/scale_ca
      -- 
    scale_ca_2669_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_0_scale_ack_1, ack => cp_elements(406)); -- 
    -- CP-element group 407 transition  output  bypass 
    -- predecessors 393 
    -- successors 408 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_883_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_883_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_883_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_1/index_resize_req
      -- 
    cp_elements(407) <= cp_elements(393);
    index_resize_req_2678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(407), ack => array_obj_ref_884_index_1_resize_req_0); -- 
    -- CP-element group 408 transition  input  output  no-bypass 
    -- predecessors 407 
    -- successors 409 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_1_resize_ack_0, ack => cp_elements(408)); -- 
    scale_rename_req_2683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(408), ack => array_obj_ref_884_index_1_rename_req_0); -- 
    -- CP-element group 409 transition  input  no-bypass 
    -- predecessors 408 
    -- successors 402 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_1_rename_ack_0, ack => cp_elements(409)); -- 
    -- CP-element group 410 transition  input  output  no-bypass 
    -- predecessors 402 
    -- successors 411 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_2689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_sum_1_ack_0, ack => cp_elements(410)); -- 
    partial_sum_1_cr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(410), ack => array_obj_ref_884_index_sum_1_req_1); -- 
    -- CP-element group 411 transition  input  output  no-bypass 
    -- predecessors 410 
    -- successors 412 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_sum_1_ack_1, ack => cp_elements(411)); -- 
    final_index_req_2692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => array_obj_ref_884_offset_inst_req_0); -- 
    -- CP-element group 412 transition  input  output  no-bypass 
    -- predecessors 411 
    -- successors 413 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_2693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_offset_inst_ack_0, ack => cp_elements(412)); -- 
    sum_rename_req_2697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(412), ack => array_obj_ref_884_root_address_inst_req_0); -- 
    -- CP-element group 413 transition  input  no-bypass 
    -- predecessors 412 
    -- successors 400 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_884_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_root_address_inst_ack_0, ack => cp_elements(413)); -- 
    -- CP-element group 414 transition  output  bypass 
    -- predecessors 400 
    -- successors 415 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_885_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_885_complete/final_reg_req
      -- 
    cp_elements(414) <= cp_elements(400);
    final_reg_req_2702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(414), ack => addr_of_885_final_reg_req_0); -- 
    -- CP-element group 415 transition  input  no-bypass 
    -- predecessors 414 
    -- successors 401 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_885_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_885_complete/final_reg_ack
      -- 
    final_reg_ack_2703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_885_final_reg_ack_0, ack => cp_elements(415)); -- 
    -- CP-element group 416 join  fork  transition  no-bypass 
    -- predecessors 418 420 
    -- successors 417 421 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_active_
      -- 
    cpelement_group_416 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(418);
      predecessors(1) <= cp_elements(420);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(416)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(416),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 417 join  fork  transition  no-bypass 
    -- predecessors 416 422 
    -- successors 431 482 557 625 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_892_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_892_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_892_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_completed_
      -- 
    cpelement_group_417 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(416);
      predecessors(1) <= cp_elements(422);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(417)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(417),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 418 fork  transition  bypass 
    -- predecessors 369 
    -- successors 416 419 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_888_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_888_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_888_completed_
      -- 
    cp_elements(418) <= cp_elements(369);
    -- CP-element group 419 transition  output  bypass 
    -- predecessors 418 
    -- successors 420 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Sample/rr
      -- 
    cp_elements(419) <= cp_elements(418);
    rr_2716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(419), ack => binary_891_inst_req_0); -- 
    -- CP-element group 420 transition  input  no-bypass 
    -- predecessors 419 
    -- successors 416 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Sample/ra
      -- 
    ra_2717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_891_inst_ack_0, ack => cp_elements(420)); -- 
    -- CP-element group 421 transition  output  bypass 
    -- predecessors 416 
    -- successors 422 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Update/cr
      -- 
    cp_elements(421) <= cp_elements(416);
    cr_2721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(421), ack => binary_891_inst_req_1); -- 
    -- CP-element group 422 transition  input  no-bypass 
    -- predecessors 421 
    -- successors 417 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_891_complete_Update/ca
      -- 
    ca_2722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_891_inst_ack_1, ack => cp_elements(422)); -- 
    -- CP-element group 423 transition  bypass 
    -- predecessors 367 
    -- successors 424 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_897_trigger_
      -- 
    cp_elements(423) <= cp_elements(367);
    -- CP-element group 424 join  fork  transition  no-bypass 
    -- predecessors 423 437 
    -- successors 425 438 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_897_active_
      -- 
    cpelement_group_424 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(423);
      predecessors(1) <= cp_elements(437);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(424)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(424),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 425 join  transition  output  bypass 
    -- predecessors 424 439 
    -- successors 1010 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_898_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_898_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_898_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_897_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1120_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1120_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1120_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_addr_resize/base_resize_req
      -- 
    cpelement_group_425 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(424);
      predecessors(1) <= cp_elements(439);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(425)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(425),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4842_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(425), ack => ptr_deref_1121_base_resize_req_0); -- 
    -- CP-element group 426 join  transition  output  bypass 
    -- predecessors 430 433 
    -- successors 434 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_426 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(430);
      predecessors(1) <= cp_elements(433);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(426)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(426),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(426), ack => array_obj_ref_896_index_sum_1_req_0); -- 
    -- CP-element group 427 transition  output  bypass 
    -- predecessors 367 
    -- successors 428 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_894_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_894_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_894_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_0/index_resize_req
      -- 
    cp_elements(427) <= cp_elements(367);
    index_resize_req_2740_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(427), ack => array_obj_ref_896_index_0_resize_req_0); -- 
    -- CP-element group 428 transition  input  output  no-bypass 
    -- predecessors 427 
    -- successors 429 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_0/scale_rr
      -- 
    index_resize_ack_2741_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_index_0_resize_ack_0, ack => cp_elements(428)); -- 
    scale_rr_2745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(428), ack => array_obj_ref_896_index_0_scale_req_0); -- 
    -- CP-element group 429 transition  input  output  no-bypass 
    -- predecessors 428 
    -- successors 430 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_0/scale_cr
      -- 
    scale_ra_2746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_index_0_scale_ack_0, ack => cp_elements(429)); -- 
    scale_cr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(429), ack => array_obj_ref_896_index_0_scale_req_1); -- 
    -- CP-element group 430 transition  input  no-bypass 
    -- predecessors 429 
    -- successors 426 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_0/scale_ca
      -- 
    scale_ca_2748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_index_0_scale_ack_1, ack => cp_elements(430)); -- 
    -- CP-element group 431 transition  output  bypass 
    -- predecessors 417 
    -- successors 432 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_895_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_895_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_895_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_1/index_resize_req
      -- 
    cp_elements(431) <= cp_elements(417);
    index_resize_req_2757_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(431), ack => array_obj_ref_896_index_1_resize_req_0); -- 
    -- CP-element group 432 transition  input  output  no-bypass 
    -- predecessors 431 
    -- successors 433 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2758_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_index_1_resize_ack_0, ack => cp_elements(432)); -- 
    scale_rename_req_2762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(432), ack => array_obj_ref_896_index_1_rename_req_0); -- 
    -- CP-element group 433 transition  input  no-bypass 
    -- predecessors 432 
    -- successors 426 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_index_1_rename_ack_0, ack => cp_elements(433)); -- 
    -- CP-element group 434 transition  input  output  no-bypass 
    -- predecessors 426 
    -- successors 435 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_2768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_index_sum_1_ack_0, ack => cp_elements(434)); -- 
    partial_sum_1_cr_2769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(434), ack => array_obj_ref_896_index_sum_1_req_1); -- 
    -- CP-element group 435 transition  input  output  no-bypass 
    -- predecessors 434 
    -- successors 436 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_index_sum_1_ack_1, ack => cp_elements(435)); -- 
    final_index_req_2771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(435), ack => array_obj_ref_896_offset_inst_req_0); -- 
    -- CP-element group 436 transition  input  output  no-bypass 
    -- predecessors 435 
    -- successors 437 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_2772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_offset_inst_ack_0, ack => cp_elements(436)); -- 
    sum_rename_req_2776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(436), ack => array_obj_ref_896_root_address_inst_req_0); -- 
    -- CP-element group 437 transition  input  no-bypass 
    -- predecessors 436 
    -- successors 424 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_896_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_896_root_address_inst_ack_0, ack => cp_elements(437)); -- 
    -- CP-element group 438 transition  output  bypass 
    -- predecessors 424 
    -- successors 439 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_897_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_897_complete/final_reg_req
      -- 
    cp_elements(438) <= cp_elements(424);
    final_reg_req_2781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(438), ack => addr_of_897_final_reg_req_0); -- 
    -- CP-element group 439 transition  input  no-bypass 
    -- predecessors 438 
    -- successors 425 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_897_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_897_complete/final_reg_ack
      -- 
    final_reg_ack_2782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_897_final_reg_ack_0, ack => cp_elements(439)); -- 
    -- CP-element group 440 transition  bypass 
    -- predecessors 367 
    -- successors 441 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_903_trigger_
      -- 
    cp_elements(440) <= cp_elements(367);
    -- CP-element group 441 join  fork  transition  no-bypass 
    -- predecessors 440 454 
    -- successors 442 455 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_903_active_
      -- 
    cpelement_group_441 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(440);
      predecessors(1) <= cp_elements(454);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(441)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(441),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 442 join  transition  output  bypass 
    -- predecessors 441 456 
    -- successors 2030 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_904_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_904_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_904_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_903_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1696_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1696_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1696_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_addr_resize/base_resize_req
      -- 
    cpelement_group_442 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(441);
      predecessors(1) <= cp_elements(456);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(442)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(442),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_8202_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(442), ack => ptr_deref_1697_base_resize_req_0); -- 
    -- CP-element group 443 join  transition  output  bypass 
    -- predecessors 447 450 
    -- successors 451 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_443 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(447);
      predecessors(1) <= cp_elements(450);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(443)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(443),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(443), ack => array_obj_ref_902_index_sum_1_req_0); -- 
    -- CP-element group 444 transition  output  bypass 
    -- predecessors 367 
    -- successors 445 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_900_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_900_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_900_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_0/index_resize_req
      -- 
    cp_elements(444) <= cp_elements(367);
    index_resize_req_2800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(444), ack => array_obj_ref_902_index_0_resize_req_0); -- 
    -- CP-element group 445 transition  input  output  no-bypass 
    -- predecessors 444 
    -- successors 446 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_0/scale_rr
      -- 
    index_resize_ack_2801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_index_0_resize_ack_0, ack => cp_elements(445)); -- 
    scale_rr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(445), ack => array_obj_ref_902_index_0_scale_req_0); -- 
    -- CP-element group 446 transition  input  output  no-bypass 
    -- predecessors 445 
    -- successors 447 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_0/scale_cr
      -- 
    scale_ra_2806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_index_0_scale_ack_0, ack => cp_elements(446)); -- 
    scale_cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(446), ack => array_obj_ref_902_index_0_scale_req_1); -- 
    -- CP-element group 447 transition  input  no-bypass 
    -- predecessors 446 
    -- successors 443 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_0/scale_ca
      -- 
    scale_ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_index_0_scale_ack_1, ack => cp_elements(447)); -- 
    -- CP-element group 448 transition  output  bypass 
    -- predecessors 369 
    -- successors 449 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_901_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_901_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_901_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_1/index_resize_req
      -- 
    cp_elements(448) <= cp_elements(369);
    index_resize_req_2817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(448), ack => array_obj_ref_902_index_1_resize_req_0); -- 
    -- CP-element group 449 transition  input  output  no-bypass 
    -- predecessors 448 
    -- successors 450 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_index_1_resize_ack_0, ack => cp_elements(449)); -- 
    scale_rename_req_2822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(449), ack => array_obj_ref_902_index_1_rename_req_0); -- 
    -- CP-element group 450 transition  input  no-bypass 
    -- predecessors 449 
    -- successors 443 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_index_1_rename_ack_0, ack => cp_elements(450)); -- 
    -- CP-element group 451 transition  input  output  no-bypass 
    -- predecessors 443 
    -- successors 452 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_2828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_index_sum_1_ack_0, ack => cp_elements(451)); -- 
    partial_sum_1_cr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(451), ack => array_obj_ref_902_index_sum_1_req_1); -- 
    -- CP-element group 452 transition  input  output  no-bypass 
    -- predecessors 451 
    -- successors 453 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_index_sum_1_ack_1, ack => cp_elements(452)); -- 
    final_index_req_2831_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(452), ack => array_obj_ref_902_offset_inst_req_0); -- 
    -- CP-element group 453 transition  input  output  no-bypass 
    -- predecessors 452 
    -- successors 454 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_2832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_offset_inst_ack_0, ack => cp_elements(453)); -- 
    sum_rename_req_2836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(453), ack => array_obj_ref_902_root_address_inst_req_0); -- 
    -- CP-element group 454 transition  input  no-bypass 
    -- predecessors 453 
    -- successors 441 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_902_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_902_root_address_inst_ack_0, ack => cp_elements(454)); -- 
    -- CP-element group 455 transition  output  bypass 
    -- predecessors 441 
    -- successors 456 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_903_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_903_complete/final_reg_req
      -- 
    cp_elements(455) <= cp_elements(441);
    final_reg_req_2841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(455), ack => addr_of_903_final_reg_req_0); -- 
    -- CP-element group 456 transition  input  no-bypass 
    -- predecessors 455 
    -- successors 442 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_903_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_903_complete/final_reg_ack
      -- 
    final_reg_ack_2842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_903_final_reg_ack_0, ack => cp_elements(456)); -- 
    -- CP-element group 457 transition  bypass 
    -- predecessors 367 
    -- successors 458 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_909_trigger_
      -- 
    cp_elements(457) <= cp_elements(367);
    -- CP-element group 458 join  fork  transition  no-bypass 
    -- predecessors 457 471 
    -- successors 459 472 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_909_active_
      -- 
    cpelement_group_458 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(457);
      predecessors(1) <= cp_elements(471);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(458)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(458),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 459 join  transition  output  bypass 
    -- predecessors 458 473 
    -- successors 2060 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_910_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_910_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_910_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_909_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1708_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1708_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1708_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_addr_resize/base_resize_req
      -- 
    cpelement_group_459 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(458);
      predecessors(1) <= cp_elements(473);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(459)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(459),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_8358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(459), ack => ptr_deref_1709_base_resize_req_0); -- 
    -- CP-element group 460 join  transition  output  bypass 
    -- predecessors 464 467 
    -- successors 468 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_460 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(464);
      predecessors(1) <= cp_elements(467);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(460)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(460),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2887_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(460), ack => array_obj_ref_908_index_sum_1_req_0); -- 
    -- CP-element group 461 transition  output  bypass 
    -- predecessors 367 
    -- successors 462 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_906_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_906_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_906_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_0/index_resize_req
      -- 
    cp_elements(461) <= cp_elements(367);
    index_resize_req_2860_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(461), ack => array_obj_ref_908_index_0_resize_req_0); -- 
    -- CP-element group 462 transition  input  output  no-bypass 
    -- predecessors 461 
    -- successors 463 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_0/scale_rr
      -- 
    index_resize_ack_2861_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_index_0_resize_ack_0, ack => cp_elements(462)); -- 
    scale_rr_2865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(462), ack => array_obj_ref_908_index_0_scale_req_0); -- 
    -- CP-element group 463 transition  input  output  no-bypass 
    -- predecessors 462 
    -- successors 464 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_0/scale_cr
      -- 
    scale_ra_2866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_index_0_scale_ack_0, ack => cp_elements(463)); -- 
    scale_cr_2867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(463), ack => array_obj_ref_908_index_0_scale_req_1); -- 
    -- CP-element group 464 transition  input  no-bypass 
    -- predecessors 463 
    -- successors 460 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_0/scale_ca
      -- 
    scale_ca_2868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_index_0_scale_ack_1, ack => cp_elements(464)); -- 
    -- CP-element group 465 transition  output  bypass 
    -- predecessors 393 
    -- successors 466 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_907_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_907_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_907_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_1/index_resize_req
      -- 
    cp_elements(465) <= cp_elements(393);
    index_resize_req_2877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(465), ack => array_obj_ref_908_index_1_resize_req_0); -- 
    -- CP-element group 466 transition  input  output  no-bypass 
    -- predecessors 465 
    -- successors 467 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_index_1_resize_ack_0, ack => cp_elements(466)); -- 
    scale_rename_req_2882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(466), ack => array_obj_ref_908_index_1_rename_req_0); -- 
    -- CP-element group 467 transition  input  no-bypass 
    -- predecessors 466 
    -- successors 460 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2883_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_index_1_rename_ack_0, ack => cp_elements(467)); -- 
    -- CP-element group 468 transition  input  output  no-bypass 
    -- predecessors 460 
    -- successors 469 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_2888_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_index_sum_1_ack_0, ack => cp_elements(468)); -- 
    partial_sum_1_cr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(468), ack => array_obj_ref_908_index_sum_1_req_1); -- 
    -- CP-element group 469 transition  input  output  no-bypass 
    -- predecessors 468 
    -- successors 470 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_index_sum_1_ack_1, ack => cp_elements(469)); -- 
    final_index_req_2891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(469), ack => array_obj_ref_908_offset_inst_req_0); -- 
    -- CP-element group 470 transition  input  output  no-bypass 
    -- predecessors 469 
    -- successors 471 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_2892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_offset_inst_ack_0, ack => cp_elements(470)); -- 
    sum_rename_req_2896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(470), ack => array_obj_ref_908_root_address_inst_req_0); -- 
    -- CP-element group 471 transition  input  no-bypass 
    -- predecessors 470 
    -- successors 458 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_908_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_908_root_address_inst_ack_0, ack => cp_elements(471)); -- 
    -- CP-element group 472 transition  output  bypass 
    -- predecessors 458 
    -- successors 473 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_909_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_909_complete/final_reg_req
      -- 
    cp_elements(472) <= cp_elements(458);
    final_reg_req_2901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(472), ack => addr_of_909_final_reg_req_0); -- 
    -- CP-element group 473 transition  input  no-bypass 
    -- predecessors 472 
    -- successors 459 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_909_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_909_complete/final_reg_ack
      -- 
    final_reg_ack_2902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_909_final_reg_ack_0, ack => cp_elements(473)); -- 
    -- CP-element group 474 transition  bypass 
    -- predecessors 367 
    -- successors 475 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_915_trigger_
      -- 
    cp_elements(474) <= cp_elements(367);
    -- CP-element group 475 join  fork  transition  no-bypass 
    -- predecessors 474 488 
    -- successors 476 489 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_915_active_
      -- 
    cpelement_group_475 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(474);
      predecessors(1) <= cp_elements(488);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(475)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(475),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 476 join  transition  output  bypass 
    -- predecessors 475 490 
    -- successors 2050 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_916_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_916_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_916_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_915_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1704_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1704_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1704_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_addr_resize/base_resize_req
      -- 
    cpelement_group_476 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(475);
      predecessors(1) <= cp_elements(490);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(476)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(476),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_8306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(476), ack => ptr_deref_1705_base_resize_req_0); -- 
    -- CP-element group 477 join  transition  output  bypass 
    -- predecessors 481 484 
    -- successors 485 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_477 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(481);
      predecessors(1) <= cp_elements(484);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(477)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(477),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_2947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(477), ack => array_obj_ref_914_index_sum_1_req_0); -- 
    -- CP-element group 478 transition  output  bypass 
    -- predecessors 367 
    -- successors 479 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_912_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_912_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_912_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_0/index_resize_req
      -- 
    cp_elements(478) <= cp_elements(367);
    index_resize_req_2920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(478), ack => array_obj_ref_914_index_0_resize_req_0); -- 
    -- CP-element group 479 transition  input  output  no-bypass 
    -- predecessors 478 
    -- successors 480 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_0/scale_rr
      -- 
    index_resize_ack_2921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_0_resize_ack_0, ack => cp_elements(479)); -- 
    scale_rr_2925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(479), ack => array_obj_ref_914_index_0_scale_req_0); -- 
    -- CP-element group 480 transition  input  output  no-bypass 
    -- predecessors 479 
    -- successors 481 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_0/scale_cr
      -- 
    scale_ra_2926_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_0_scale_ack_0, ack => cp_elements(480)); -- 
    scale_cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(480), ack => array_obj_ref_914_index_0_scale_req_1); -- 
    -- CP-element group 481 transition  input  no-bypass 
    -- predecessors 480 
    -- successors 477 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_0/scale_ca
      -- 
    scale_ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_0_scale_ack_1, ack => cp_elements(481)); -- 
    -- CP-element group 482 transition  output  bypass 
    -- predecessors 417 
    -- successors 483 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_913_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_913_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_913_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_1/index_resize_req
      -- 
    cp_elements(482) <= cp_elements(417);
    index_resize_req_2937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(482), ack => array_obj_ref_914_index_1_resize_req_0); -- 
    -- CP-element group 483 transition  input  output  no-bypass 
    -- predecessors 482 
    -- successors 484 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_2938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_1_resize_ack_0, ack => cp_elements(483)); -- 
    scale_rename_req_2942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(483), ack => array_obj_ref_914_index_1_rename_req_0); -- 
    -- CP-element group 484 transition  input  no-bypass 
    -- predecessors 483 
    -- successors 477 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_2943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_1_rename_ack_0, ack => cp_elements(484)); -- 
    -- CP-element group 485 transition  input  output  no-bypass 
    -- predecessors 477 
    -- successors 486 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_2948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_sum_1_ack_0, ack => cp_elements(485)); -- 
    partial_sum_1_cr_2949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(485), ack => array_obj_ref_914_index_sum_1_req_1); -- 
    -- CP-element group 486 transition  input  output  no-bypass 
    -- predecessors 485 
    -- successors 487 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/final_index_req
      -- 
    partial_sum_1_ca_2950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_index_sum_1_ack_1, ack => cp_elements(486)); -- 
    final_index_req_2951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(486), ack => array_obj_ref_914_offset_inst_req_0); -- 
    -- CP-element group 487 transition  input  output  no-bypass 
    -- predecessors 486 
    -- successors 488 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_2952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_offset_inst_ack_0, ack => cp_elements(487)); -- 
    sum_rename_req_2956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(487), ack => array_obj_ref_914_root_address_inst_req_0); -- 
    -- CP-element group 488 transition  input  no-bypass 
    -- predecessors 487 
    -- successors 475 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_914_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_914_root_address_inst_ack_0, ack => cp_elements(488)); -- 
    -- CP-element group 489 transition  output  bypass 
    -- predecessors 475 
    -- successors 490 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_915_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_915_complete/$entry
      -- 
    cp_elements(489) <= cp_elements(475);
    final_reg_req_2961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(489), ack => addr_of_915_final_reg_req_0); -- 
    -- CP-element group 490 transition  input  no-bypass 
    -- predecessors 489 
    -- successors 476 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_915_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_915_complete/$exit
      -- 
    final_reg_ack_2962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_915_final_reg_ack_0, ack => cp_elements(490)); -- 
    -- CP-element group 491 join  fork  transition  no-bypass 
    -- predecessors 493 495 
    -- successors 492 496 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_active_
      -- 
    cpelement_group_491 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(493);
      predecessors(1) <= cp_elements(495);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(491)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(491),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 492 join  fork  transition  no-bypass 
    -- predecessors 491 497 
    -- successors 506 574 642 659 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_922_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_922_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_922_trigger_
      -- 
    cpelement_group_492 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(491);
      predecessors(1) <= cp_elements(497);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(492)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(492),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 493 fork  transition  bypass 
    -- predecessors 369 
    -- successors 491 494 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_918_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_918_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_918_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_trigger_
      -- 
    cp_elements(493) <= cp_elements(369);
    -- CP-element group 494 transition  output  bypass 
    -- predecessors 493 
    -- successors 495 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Sample/$entry
      -- 
    cp_elements(494) <= cp_elements(493);
    rr_2975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(494), ack => binary_921_inst_req_0); -- 
    -- CP-element group 495 transition  input  no-bypass 
    -- predecessors 494 
    -- successors 491 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Sample/$exit
      -- 
    ra_2976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_921_inst_ack_0, ack => cp_elements(495)); -- 
    -- CP-element group 496 transition  output  bypass 
    -- predecessors 491 
    -- successors 497 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Update/$entry
      -- 
    cp_elements(496) <= cp_elements(491);
    cr_2980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(496), ack => binary_921_inst_req_1); -- 
    -- CP-element group 497 transition  input  no-bypass 
    -- predecessors 496 
    -- successors 492 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_921_complete_Update/$exit
      -- 
    ca_2981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_921_inst_ack_1, ack => cp_elements(497)); -- 
    -- CP-element group 498 transition  bypass 
    -- predecessors 367 
    -- successors 499 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_927_trigger_
      -- 
    cp_elements(498) <= cp_elements(367);
    -- CP-element group 499 join  fork  transition  no-bypass 
    -- predecessors 498 512 
    -- successors 500 513 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_927_active_
      -- 
    cpelement_group_499 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(498);
      predecessors(1) <= cp_elements(512);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(499)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(499),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 500 join  transition  output  bypass 
    -- predecessors 499 514 
    -- successors 2040 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_927_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_928_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_928_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_928_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1700_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1700_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1700_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_addr_resize/base_resize_req
      -- 
    cpelement_group_500 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(499);
      predecessors(1) <= cp_elements(514);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(500)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(500),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_8254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => ptr_deref_1701_base_resize_req_0); -- 
    -- CP-element group 501 join  transition  output  bypass 
    -- predecessors 505 508 
    -- successors 509 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_indices_scaled
      -- 
    cpelement_group_501 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(505);
      predecessors(1) <= cp_elements(508);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(501)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(501),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(501), ack => array_obj_ref_926_index_sum_1_req_0); -- 
    -- CP-element group 502 transition  output  bypass 
    -- predecessors 367 
    -- successors 503 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_924_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_924_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_924_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_computed_0
      -- 
    cp_elements(502) <= cp_elements(367);
    index_resize_req_2999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(502), ack => array_obj_ref_926_index_0_resize_req_0); -- 
    -- CP-element group 503 transition  input  output  no-bypass 
    -- predecessors 502 
    -- successors 504 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resized_0
      -- 
    index_resize_ack_3000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_index_0_resize_ack_0, ack => cp_elements(503)); -- 
    scale_rr_3004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(503), ack => array_obj_ref_926_index_0_scale_req_0); -- 
    -- CP-element group 504 transition  input  output  no-bypass 
    -- predecessors 503 
    -- successors 505 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_0/scale_ra
      -- 
    scale_ra_3005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_index_0_scale_ack_0, ack => cp_elements(504)); -- 
    scale_cr_3006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(504), ack => array_obj_ref_926_index_0_scale_req_1); -- 
    -- CP-element group 505 transition  input  no-bypass 
    -- predecessors 504 
    -- successors 501 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_0/$exit
      -- 
    scale_ca_3007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_index_0_scale_ack_1, ack => cp_elements(505)); -- 
    -- CP-element group 506 transition  output  bypass 
    -- predecessors 492 
    -- successors 507 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_925_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_925_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_925_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_computed_1
      -- 
    cp_elements(506) <= cp_elements(492);
    index_resize_req_3016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => array_obj_ref_926_index_1_resize_req_0); -- 
    -- CP-element group 507 transition  input  output  no-bypass 
    -- predecessors 506 
    -- successors 508 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_resized_1
      -- 
    index_resize_ack_3017_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_index_1_resize_ack_0, ack => cp_elements(507)); -- 
    scale_rename_req_3021_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(507), ack => array_obj_ref_926_index_1_rename_req_0); -- 
    -- CP-element group 508 transition  input  no-bypass 
    -- predecessors 507 
    -- successors 501 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_index_scale_1/$exit
      -- 
    scale_rename_ack_3022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_index_1_rename_ack_0, ack => cp_elements(508)); -- 
    -- CP-element group 509 transition  input  output  no-bypass 
    -- predecessors 501 
    -- successors 510 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_3027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_index_sum_1_ack_0, ack => cp_elements(509)); -- 
    partial_sum_1_cr_3028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => array_obj_ref_926_index_sum_1_req_1); -- 
    -- CP-element group 510 transition  input  output  no-bypass 
    -- predecessors 509 
    -- successors 511 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_3029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_index_sum_1_ack_1, ack => cp_elements(510)); -- 
    final_index_req_3030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(510), ack => array_obj_ref_926_offset_inst_req_0); -- 
    -- CP-element group 511 transition  input  output  no-bypass 
    -- predecessors 510 
    -- successors 512 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_offset_calculated
      -- 
    final_index_ack_3031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_offset_inst_ack_0, ack => cp_elements(511)); -- 
    sum_rename_req_3035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(511), ack => array_obj_ref_926_root_address_inst_req_0); -- 
    -- CP-element group 512 transition  input  no-bypass 
    -- predecessors 511 
    -- successors 499 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_926_root_address_calculated
      -- 
    sum_rename_ack_3036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_926_root_address_inst_ack_0, ack => cp_elements(512)); -- 
    -- CP-element group 513 transition  output  bypass 
    -- predecessors 499 
    -- successors 514 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_927_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_927_complete/$entry
      -- 
    cp_elements(513) <= cp_elements(499);
    final_reg_req_3040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(513), ack => addr_of_927_final_reg_req_0); -- 
    -- CP-element group 514 transition  input  no-bypass 
    -- predecessors 513 
    -- successors 500 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_927_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_927_complete/$exit
      -- 
    final_reg_ack_3041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_927_final_reg_ack_0, ack => cp_elements(514)); -- 
    -- CP-element group 515 transition  bypass 
    -- predecessors 367 
    -- successors 516 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_933_trigger_
      -- 
    cp_elements(515) <= cp_elements(367);
    -- CP-element group 516 join  fork  transition  no-bypass 
    -- predecessors 515 529 
    -- successors 517 530 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_933_active_
      -- 
    cpelement_group_516 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(515);
      predecessors(1) <= cp_elements(529);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(516)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(516),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 517 join  transition  output  bypass 
    -- predecessors 516 531 
    -- successors 1730 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_933_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_934_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_934_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_934_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1520_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1520_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1520_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_addr_resize/base_resize_req
      -- 
    cpelement_group_517 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(516);
      predecessors(1) <= cp_elements(531);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(517)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(517),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_7290_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(517), ack => ptr_deref_1521_base_resize_req_0); -- 
    -- CP-element group 518 join  transition  output  bypass 
    -- predecessors 522 525 
    -- successors 526 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_indices_scaled
      -- 
    cpelement_group_518 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(522);
      predecessors(1) <= cp_elements(525);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(518)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(518),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(518), ack => array_obj_ref_932_index_sum_1_req_0); -- 
    -- CP-element group 519 transition  output  bypass 
    -- predecessors 367 
    -- successors 520 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_930_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_930_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_930_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_computed_0
      -- 
    cp_elements(519) <= cp_elements(367);
    index_resize_req_3059_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(519), ack => array_obj_ref_932_index_0_resize_req_0); -- 
    -- CP-element group 520 transition  input  output  no-bypass 
    -- predecessors 519 
    -- successors 521 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resized_0
      -- 
    index_resize_ack_3060_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_0_resize_ack_0, ack => cp_elements(520)); -- 
    scale_rr_3064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(520), ack => array_obj_ref_932_index_0_scale_req_0); -- 
    -- CP-element group 521 transition  input  output  no-bypass 
    -- predecessors 520 
    -- successors 522 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_0/scale_ra
      -- 
    scale_ra_3065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_0_scale_ack_0, ack => cp_elements(521)); -- 
    scale_cr_3066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(521), ack => array_obj_ref_932_index_0_scale_req_1); -- 
    -- CP-element group 522 transition  input  no-bypass 
    -- predecessors 521 
    -- successors 518 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_0/$exit
      -- 
    scale_ca_3067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_0_scale_ack_1, ack => cp_elements(522)); -- 
    -- CP-element group 523 transition  output  bypass 
    -- predecessors 369 
    -- successors 524 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_931_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_931_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_931_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_1/index_resize_req
      -- 
    cp_elements(523) <= cp_elements(369);
    index_resize_req_3076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(523), ack => array_obj_ref_932_index_1_resize_req_0); -- 
    -- CP-element group 524 transition  input  output  no-bypass 
    -- predecessors 523 
    -- successors 525 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_1_resize_ack_0, ack => cp_elements(524)); -- 
    scale_rename_req_3081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(524), ack => array_obj_ref_932_index_1_rename_req_0); -- 
    -- CP-element group 525 transition  input  no-bypass 
    -- predecessors 524 
    -- successors 518 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_index_scale_1/$exit
      -- 
    scale_rename_ack_3082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_1_rename_ack_0, ack => cp_elements(525)); -- 
    -- CP-element group 526 transition  input  output  no-bypass 
    -- predecessors 518 
    -- successors 527 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_sum_1_ack_0, ack => cp_elements(526)); -- 
    partial_sum_1_cr_3088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(526), ack => array_obj_ref_932_index_sum_1_req_1); -- 
    -- CP-element group 527 transition  input  output  no-bypass 
    -- predecessors 526 
    -- successors 528 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_3089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_sum_1_ack_1, ack => cp_elements(527)); -- 
    final_index_req_3090_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(527), ack => array_obj_ref_932_offset_inst_req_0); -- 
    -- CP-element group 528 transition  input  output  no-bypass 
    -- predecessors 527 
    -- successors 529 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_offset_calculated
      -- 
    final_index_ack_3091_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_offset_inst_ack_0, ack => cp_elements(528)); -- 
    sum_rename_req_3095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(528), ack => array_obj_ref_932_root_address_inst_req_0); -- 
    -- CP-element group 529 transition  input  no-bypass 
    -- predecessors 528 
    -- successors 516 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_932_root_address_calculated
      -- 
    sum_rename_ack_3096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_root_address_inst_ack_0, ack => cp_elements(529)); -- 
    -- CP-element group 530 transition  output  bypass 
    -- predecessors 516 
    -- successors 531 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_933_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_933_complete/$entry
      -- 
    cp_elements(530) <= cp_elements(516);
    final_reg_req_3100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(530), ack => addr_of_933_final_reg_req_0); -- 
    -- CP-element group 531 transition  input  no-bypass 
    -- predecessors 530 
    -- successors 517 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_933_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_933_complete/$exit
      -- 
    final_reg_ack_3101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_933_final_reg_ack_0, ack => cp_elements(531)); -- 
    -- CP-element group 532 transition  bypass 
    -- predecessors 367 
    -- successors 533 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_939_trigger_
      -- 
    cp_elements(532) <= cp_elements(367);
    -- CP-element group 533 join  fork  transition  no-bypass 
    -- predecessors 532 546 
    -- successors 534 547 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_939_active_
      -- 
    cpelement_group_533 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(532);
      predecessors(1) <= cp_elements(546);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(533)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(533),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 534 join  transition  output  bypass 
    -- predecessors 533 548 
    -- successors 1760 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_940_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_940_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_940_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_939_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1532_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1532_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1532_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_addr_resize/base_resize_req
      -- 
    cpelement_group_534 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(533);
      predecessors(1) <= cp_elements(548);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(534)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(534),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_7446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(534), ack => ptr_deref_1533_base_resize_req_0); -- 
    -- CP-element group 535 join  transition  output  bypass 
    -- predecessors 539 542 
    -- successors 543 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/$entry
      -- 
    cpelement_group_535 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(539);
      predecessors(1) <= cp_elements(542);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(535)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(535),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(535), ack => array_obj_ref_938_index_sum_1_req_0); -- 
    -- CP-element group 536 transition  output  bypass 
    -- predecessors 367 
    -- successors 537 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_936_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_936_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_936_completed_
      -- 
    cp_elements(536) <= cp_elements(367);
    index_resize_req_3119_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(536), ack => array_obj_ref_938_index_0_resize_req_0); -- 
    -- CP-element group 537 transition  input  output  no-bypass 
    -- predecessors 536 
    -- successors 538 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_0/$exit
      -- 
    index_resize_ack_3120_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_0_resize_ack_0, ack => cp_elements(537)); -- 
    scale_rr_3124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(537), ack => array_obj_ref_938_index_0_scale_req_0); -- 
    -- CP-element group 538 transition  input  output  no-bypass 
    -- predecessors 537 
    -- successors 539 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_0/scale_ra
      -- 
    scale_ra_3125_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_0_scale_ack_0, ack => cp_elements(538)); -- 
    scale_cr_3126_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(538), ack => array_obj_ref_938_index_0_scale_req_1); -- 
    -- CP-element group 539 transition  input  no-bypass 
    -- predecessors 538 
    -- successors 535 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_0/$exit
      -- 
    scale_ca_3127_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_0_scale_ack_1, ack => cp_elements(539)); -- 
    -- CP-element group 540 transition  output  bypass 
    -- predecessors 393 
    -- successors 541 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_937_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_937_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_937_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_computed_1
      -- 
    cp_elements(540) <= cp_elements(393);
    index_resize_req_3136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(540), ack => array_obj_ref_938_index_1_resize_req_0); -- 
    -- CP-element group 541 transition  input  output  no-bypass 
    -- predecessors 540 
    -- successors 542 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_resized_1
      -- 
    index_resize_ack_3137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_1_resize_ack_0, ack => cp_elements(541)); -- 
    scale_rename_req_3141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => array_obj_ref_938_index_1_rename_req_0); -- 
    -- CP-element group 542 transition  input  no-bypass 
    -- predecessors 541 
    -- successors 535 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_index_scale_1/$exit
      -- 
    scale_rename_ack_3142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_1_rename_ack_0, ack => cp_elements(542)); -- 
    -- CP-element group 543 transition  input  output  no-bypass 
    -- predecessors 535 
    -- successors 544 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_3147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_sum_1_ack_0, ack => cp_elements(543)); -- 
    partial_sum_1_cr_3148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(543), ack => array_obj_ref_938_index_sum_1_req_1); -- 
    -- CP-element group 544 transition  input  output  no-bypass 
    -- predecessors 543 
    -- successors 545 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_3149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_index_sum_1_ack_1, ack => cp_elements(544)); -- 
    final_index_req_3150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(544), ack => array_obj_ref_938_offset_inst_req_0); -- 
    -- CP-element group 545 transition  input  output  no-bypass 
    -- predecessors 544 
    -- successors 546 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_add_indices/$exit
      -- 
    final_index_ack_3151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_offset_inst_ack_0, ack => cp_elements(545)); -- 
    sum_rename_req_3155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(545), ack => array_obj_ref_938_root_address_inst_req_0); -- 
    -- CP-element group 546 transition  input  no-bypass 
    -- predecessors 545 
    -- successors 533 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_938_base_plus_offset/$exit
      -- 
    sum_rename_ack_3156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_938_root_address_inst_ack_0, ack => cp_elements(546)); -- 
    -- CP-element group 547 transition  output  bypass 
    -- predecessors 533 
    -- successors 548 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_939_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_939_complete/$entry
      -- 
    cp_elements(547) <= cp_elements(533);
    final_reg_req_3160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(547), ack => addr_of_939_final_reg_req_0); -- 
    -- CP-element group 548 transition  input  no-bypass 
    -- predecessors 547 
    -- successors 534 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_939_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_939_complete/$exit
      -- 
    final_reg_ack_3161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_939_final_reg_ack_0, ack => cp_elements(548)); -- 
    -- CP-element group 549 transition  bypass 
    -- predecessors 367 
    -- successors 550 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_945_trigger_
      -- 
    cp_elements(549) <= cp_elements(367);
    -- CP-element group 550 join  fork  transition  no-bypass 
    -- predecessors 549 563 
    -- successors 551 564 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_945_active_
      -- 
    cpelement_group_550 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(549);
      predecessors(1) <= cp_elements(563);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(550)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(550),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 551 join  transition  output  bypass 
    -- predecessors 550 565 
    -- successors 1750 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_945_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_946_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_946_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_946_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1528_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1528_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1528_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_addr_resize/base_resize_req
      -- 
    cpelement_group_551 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(550);
      predecessors(1) <= cp_elements(565);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(551)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(551),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_7394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(551), ack => ptr_deref_1529_base_resize_req_0); -- 
    -- CP-element group 552 join  transition  output  bypass 
    -- predecessors 556 559 
    -- successors 560 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/$entry
      -- 
    cpelement_group_552 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(556);
      predecessors(1) <= cp_elements(559);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(552)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(552),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3206_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(552), ack => array_obj_ref_944_index_sum_1_req_0); -- 
    -- CP-element group 553 transition  output  bypass 
    -- predecessors 367 
    -- successors 554 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_942_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_942_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_942_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_computed_0
      -- 
    cp_elements(553) <= cp_elements(367);
    index_resize_req_3179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(553), ack => array_obj_ref_944_index_0_resize_req_0); -- 
    -- CP-element group 554 transition  input  output  no-bypass 
    -- predecessors 553 
    -- successors 555 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resized_0
      -- 
    index_resize_ack_3180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_index_0_resize_ack_0, ack => cp_elements(554)); -- 
    scale_rr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(554), ack => array_obj_ref_944_index_0_scale_req_0); -- 
    -- CP-element group 555 transition  input  output  no-bypass 
    -- predecessors 554 
    -- successors 556 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_0/scale_cr
      -- 
    scale_ra_3185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_index_0_scale_ack_0, ack => cp_elements(555)); -- 
    scale_cr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(555), ack => array_obj_ref_944_index_0_scale_req_1); -- 
    -- CP-element group 556 transition  input  no-bypass 
    -- predecessors 555 
    -- successors 552 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_0/scale_ca
      -- 
    scale_ca_3187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_index_0_scale_ack_1, ack => cp_elements(556)); -- 
    -- CP-element group 557 transition  output  bypass 
    -- predecessors 417 
    -- successors 558 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_943_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_943_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_943_completed_
      -- 
    cp_elements(557) <= cp_elements(417);
    index_resize_req_3196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(557), ack => array_obj_ref_944_index_1_resize_req_0); -- 
    -- CP-element group 558 transition  input  output  no-bypass 
    -- predecessors 557 
    -- successors 559 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_resize_1/$exit
      -- 
    index_resize_ack_3197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_index_1_resize_ack_0, ack => cp_elements(558)); -- 
    scale_rename_req_3201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(558), ack => array_obj_ref_944_index_1_rename_req_0); -- 
    -- CP-element group 559 transition  input  no-bypass 
    -- predecessors 558 
    -- successors 552 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_index_scale_1/$exit
      -- 
    scale_rename_ack_3202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_index_1_rename_ack_0, ack => cp_elements(559)); -- 
    -- CP-element group 560 transition  input  output  no-bypass 
    -- predecessors 552 
    -- successors 561 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_3207_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_index_sum_1_ack_0, ack => cp_elements(560)); -- 
    partial_sum_1_cr_3208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(560), ack => array_obj_ref_944_index_sum_1_req_1); -- 
    -- CP-element group 561 transition  input  output  no-bypass 
    -- predecessors 560 
    -- successors 562 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_3209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_index_sum_1_ack_1, ack => cp_elements(561)); -- 
    final_index_req_3210_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(561), ack => array_obj_ref_944_offset_inst_req_0); -- 
    -- CP-element group 562 transition  input  output  no-bypass 
    -- predecessors 561 
    -- successors 563 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_add_indices/$exit
      -- 
    final_index_ack_3211_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_offset_inst_ack_0, ack => cp_elements(562)); -- 
    sum_rename_req_3215_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(562), ack => array_obj_ref_944_root_address_inst_req_0); -- 
    -- CP-element group 563 transition  input  no-bypass 
    -- predecessors 562 
    -- successors 550 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_944_base_plus_offset/$exit
      -- 
    sum_rename_ack_3216_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_944_root_address_inst_ack_0, ack => cp_elements(563)); -- 
    -- CP-element group 564 transition  output  bypass 
    -- predecessors 550 
    -- successors 565 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_945_complete/final_reg_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_945_complete/$entry
      -- 
    cp_elements(564) <= cp_elements(550);
    final_reg_req_3220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(564), ack => addr_of_945_final_reg_req_0); -- 
    -- CP-element group 565 transition  input  no-bypass 
    -- predecessors 564 
    -- successors 551 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_945_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_945_complete/$exit
      -- 
    final_reg_ack_3221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_945_final_reg_ack_0, ack => cp_elements(565)); -- 
    -- CP-element group 566 transition  bypass 
    -- predecessors 367 
    -- successors 567 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_951_trigger_
      -- 
    cp_elements(566) <= cp_elements(367);
    -- CP-element group 567 join  fork  transition  no-bypass 
    -- predecessors 566 580 
    -- successors 568 581 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_951_active_
      -- 
    cpelement_group_567 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(566);
      predecessors(1) <= cp_elements(580);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(567)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(567),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 568 join  transition  output  bypass 
    -- predecessors 567 582 
    -- successors 1740 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_952_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_952_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_951_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_952_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1524_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1524_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1524_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_addr_resize/base_resize_req
      -- 
    cpelement_group_568 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(567);
      predecessors(1) <= cp_elements(582);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(568)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(568),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_7342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(568), ack => ptr_deref_1525_base_resize_req_0); -- 
    -- CP-element group 569 join  transition  output  bypass 
    -- predecessors 573 576 
    -- successors 577 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/$entry
      -- 
    cpelement_group_569 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(573);
      predecessors(1) <= cp_elements(576);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(569)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(569),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(569), ack => array_obj_ref_950_index_sum_1_req_0); -- 
    -- CP-element group 570 transition  output  bypass 
    -- predecessors 367 
    -- successors 571 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_948_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_948_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_948_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_0/$entry
      -- 
    cp_elements(570) <= cp_elements(367);
    index_resize_req_3239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(570), ack => array_obj_ref_950_index_0_resize_req_0); -- 
    -- CP-element group 571 transition  input  output  no-bypass 
    -- predecessors 570 
    -- successors 572 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_0/scale_rr
      -- 
    index_resize_ack_3240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_0_resize_ack_0, ack => cp_elements(571)); -- 
    scale_rr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => array_obj_ref_950_index_0_scale_req_0); -- 
    -- CP-element group 572 transition  input  output  no-bypass 
    -- predecessors 571 
    -- successors 573 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_0/scale_cr
      -- 
    scale_ra_3245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_0_scale_ack_0, ack => cp_elements(572)); -- 
    scale_cr_3246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(572), ack => array_obj_ref_950_index_0_scale_req_1); -- 
    -- CP-element group 573 transition  input  no-bypass 
    -- predecessors 572 
    -- successors 569 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_0/$exit
      -- 
    scale_ca_3247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_0_scale_ack_1, ack => cp_elements(573)); -- 
    -- CP-element group 574 transition  output  bypass 
    -- predecessors 492 
    -- successors 575 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_949_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_949_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_949_trigger_
      -- 
    cp_elements(574) <= cp_elements(492);
    index_resize_req_3256_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(574), ack => array_obj_ref_950_index_1_resize_req_0); -- 
    -- CP-element group 575 transition  input  output  no-bypass 
    -- predecessors 574 
    -- successors 576 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3257_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_1_resize_ack_0, ack => cp_elements(575)); -- 
    scale_rename_req_3261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(575), ack => array_obj_ref_950_index_1_rename_req_0); -- 
    -- CP-element group 576 transition  input  no-bypass 
    -- predecessors 575 
    -- successors 569 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_index_scale_1/$exit
      -- 
    scale_rename_ack_3262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_1_rename_ack_0, ack => cp_elements(576)); -- 
    -- CP-element group 577 transition  input  output  no-bypass 
    -- predecessors 569 
    -- successors 578 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_3267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_sum_1_ack_0, ack => cp_elements(577)); -- 
    partial_sum_1_cr_3268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(577), ack => array_obj_ref_950_index_sum_1_req_1); -- 
    -- CP-element group 578 transition  input  output  no-bypass 
    -- predecessors 577 
    -- successors 579 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/final_index_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/partial_sum_1_ca
      -- 
    partial_sum_1_ca_3269_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_index_sum_1_ack_1, ack => cp_elements(578)); -- 
    final_index_req_3270_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(578), ack => array_obj_ref_950_offset_inst_req_0); -- 
    -- CP-element group 579 transition  input  output  no-bypass 
    -- predecessors 578 
    -- successors 580 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_add_indices/$exit
      -- 
    final_index_ack_3271_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_offset_inst_ack_0, ack => cp_elements(579)); -- 
    sum_rename_req_3275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(579), ack => array_obj_ref_950_root_address_inst_req_0); -- 
    -- CP-element group 580 transition  input  no-bypass 
    -- predecessors 579 
    -- successors 567 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_950_root_address_calculated
      -- 
    sum_rename_ack_3276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_950_root_address_inst_ack_0, ack => cp_elements(580)); -- 
    -- CP-element group 581 transition  output  bypass 
    -- predecessors 567 
    -- successors 582 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_951_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_951_complete/final_reg_req
      -- 
    cp_elements(581) <= cp_elements(567);
    final_reg_req_3280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(581), ack => addr_of_951_final_reg_req_0); -- 
    -- CP-element group 582 transition  input  no-bypass 
    -- predecessors 581 
    -- successors 568 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_951_complete/final_reg_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_951_complete/$exit
      -- 
    final_reg_ack_3281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_951_final_reg_ack_0, ack => cp_elements(582)); -- 
    -- CP-element group 583 transition  bypass 
    -- predecessors 367 
    -- successors 584 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_957_trigger_
      -- 
    cp_elements(583) <= cp_elements(367);
    -- CP-element group 584 join  fork  transition  no-bypass 
    -- predecessors 583 597 
    -- successors 585 598 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_957_active_
      -- 
    cpelement_group_584 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(583);
      predecessors(1) <= cp_elements(597);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(584)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(584),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 585 join  transition  output  bypass 
    -- predecessors 584 599 
    -- successors 1430 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_958_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_957_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_958_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_958_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1344_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1344_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1344_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_addr_resize/base_resize_req
      -- 
    cpelement_group_585 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(584);
      predecessors(1) <= cp_elements(599);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(585)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(585),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_6378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(585), ack => ptr_deref_1345_base_resize_req_0); -- 
    -- CP-element group 586 join  transition  output  bypass 
    -- predecessors 590 593 
    -- successors 594 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_586 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(590);
      predecessors(1) <= cp_elements(593);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(586)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(586),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(586), ack => array_obj_ref_956_index_sum_1_req_0); -- 
    -- CP-element group 587 transition  output  bypass 
    -- predecessors 367 
    -- successors 588 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_954_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_954_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_954_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_computed_0
      -- 
    cp_elements(587) <= cp_elements(367);
    index_resize_req_3299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(587), ack => array_obj_ref_956_index_0_resize_req_0); -- 
    -- CP-element group 588 transition  input  output  no-bypass 
    -- predecessors 587 
    -- successors 589 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resized_0
      -- 
    index_resize_ack_3300_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_0_resize_ack_0, ack => cp_elements(588)); -- 
    scale_rr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(588), ack => array_obj_ref_956_index_0_scale_req_0); -- 
    -- CP-element group 589 transition  input  output  no-bypass 
    -- predecessors 588 
    -- successors 590 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_0/scale_cr
      -- 
    scale_ra_3305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_0_scale_ack_0, ack => cp_elements(589)); -- 
    scale_cr_3306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(589), ack => array_obj_ref_956_index_0_scale_req_1); -- 
    -- CP-element group 590 transition  input  no-bypass 
    -- predecessors 589 
    -- successors 586 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_0/$exit
      -- 
    scale_ca_3307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_0_scale_ack_1, ack => cp_elements(590)); -- 
    -- CP-element group 591 transition  output  bypass 
    -- predecessors 369 
    -- successors 592 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_955_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_955_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_955_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_1/$entry
      -- 
    cp_elements(591) <= cp_elements(369);
    index_resize_req_3316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => array_obj_ref_956_index_1_resize_req_0); -- 
    -- CP-element group 592 transition  input  output  no-bypass 
    -- predecessors 591 
    -- successors 593 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_resize_1/$exit
      -- 
    index_resize_ack_3317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_1_resize_ack_0, ack => cp_elements(592)); -- 
    scale_rename_req_3321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(592), ack => array_obj_ref_956_index_1_rename_req_0); -- 
    -- CP-element group 593 transition  input  no-bypass 
    -- predecessors 592 
    -- successors 586 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_index_scale_1/$exit
      -- 
    scale_rename_ack_3322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_1_rename_ack_0, ack => cp_elements(593)); -- 
    -- CP-element group 594 transition  input  output  no-bypass 
    -- predecessors 586 
    -- successors 595 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_3327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_sum_1_ack_0, ack => cp_elements(594)); -- 
    partial_sum_1_cr_3328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(594), ack => array_obj_ref_956_index_sum_1_req_1); -- 
    -- CP-element group 595 transition  input  output  no-bypass 
    -- predecessors 594 
    -- successors 596 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_index_sum_1_ack_1, ack => cp_elements(595)); -- 
    final_index_req_3330_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(595), ack => array_obj_ref_956_offset_inst_req_0); -- 
    -- CP-element group 596 transition  input  output  no-bypass 
    -- predecessors 595 
    -- successors 597 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_add_indices/$exit
      -- 
    final_index_ack_3331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_offset_inst_ack_0, ack => cp_elements(596)); -- 
    sum_rename_req_3335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(596), ack => array_obj_ref_956_root_address_inst_req_0); -- 
    -- CP-element group 597 transition  input  no-bypass 
    -- predecessors 596 
    -- successors 584 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_956_base_plus_offset/$exit
      -- 
    sum_rename_ack_3336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_956_root_address_inst_ack_0, ack => cp_elements(597)); -- 
    -- CP-element group 598 transition  output  bypass 
    -- predecessors 584 
    -- successors 599 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_957_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_957_complete/final_reg_req
      -- 
    cp_elements(598) <= cp_elements(584);
    final_reg_req_3340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(598), ack => addr_of_957_final_reg_req_0); -- 
    -- CP-element group 599 transition  input  no-bypass 
    -- predecessors 598 
    -- successors 585 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_957_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_957_complete/final_reg_ack
      -- 
    final_reg_ack_3341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_957_final_reg_ack_0, ack => cp_elements(599)); -- 
    -- CP-element group 600 transition  bypass 
    -- predecessors 367 
    -- successors 601 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_963_trigger_
      -- 
    cp_elements(600) <= cp_elements(367);
    -- CP-element group 601 join  fork  transition  no-bypass 
    -- predecessors 600 614 
    -- successors 602 615 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_963_active_
      -- 
    cpelement_group_601 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(600);
      predecessors(1) <= cp_elements(614);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(601)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(601),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 602 join  transition  output  bypass 
    -- predecessors 601 616 
    -- successors 1460 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_963_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_964_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_964_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_964_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1356_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1356_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1356_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_addr_resize/base_resize_req
      -- 
    cpelement_group_602 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(601);
      predecessors(1) <= cp_elements(616);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(602)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(602),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_6534_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(602), ack => ptr_deref_1357_base_resize_req_0); -- 
    -- CP-element group 603 join  transition  output  bypass 
    -- predecessors 607 610 
    -- successors 611 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_603 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(607);
      predecessors(1) <= cp_elements(610);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(603)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(603),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(603), ack => array_obj_ref_962_index_sum_1_req_0); -- 
    -- CP-element group 604 transition  output  bypass 
    -- predecessors 367 
    -- successors 605 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_960_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_960_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_960_completed_
      -- 
    cp_elements(604) <= cp_elements(367);
    index_resize_req_3359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(604), ack => array_obj_ref_962_index_0_resize_req_0); -- 
    -- CP-element group 605 transition  input  output  no-bypass 
    -- predecessors 604 
    -- successors 606 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_0/$entry
      -- 
    index_resize_ack_3360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_index_0_resize_ack_0, ack => cp_elements(605)); -- 
    scale_rr_3364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(605), ack => array_obj_ref_962_index_0_scale_req_0); -- 
    -- CP-element group 606 transition  input  output  no-bypass 
    -- predecessors 605 
    -- successors 607 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_0/scale_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_0/scale_ra
      -- 
    scale_ra_3365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_index_0_scale_ack_0, ack => cp_elements(606)); -- 
    scale_cr_3366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(606), ack => array_obj_ref_962_index_0_scale_req_1); -- 
    -- CP-element group 607 transition  input  no-bypass 
    -- predecessors 606 
    -- successors 603 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_0/scale_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_0/$exit
      -- 
    scale_ca_3367_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_index_0_scale_ack_1, ack => cp_elements(607)); -- 
    -- CP-element group 608 transition  output  bypass 
    -- predecessors 393 
    -- successors 609 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_961_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_961_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_961_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_1/$entry
      -- 
    cp_elements(608) <= cp_elements(393);
    index_resize_req_3376_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(608), ack => array_obj_ref_962_index_1_resize_req_0); -- 
    -- CP-element group 609 transition  input  output  no-bypass 
    -- predecessors 608 
    -- successors 610 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3377_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_index_1_resize_ack_0, ack => cp_elements(609)); -- 
    scale_rename_req_3381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(609), ack => array_obj_ref_962_index_1_rename_req_0); -- 
    -- CP-element group 610 transition  input  no-bypass 
    -- predecessors 609 
    -- successors 603 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_index_1_rename_ack_0, ack => cp_elements(610)); -- 
    -- CP-element group 611 transition  input  output  no-bypass 
    -- predecessors 603 
    -- successors 612 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_index_sum_1_ack_0, ack => cp_elements(611)); -- 
    partial_sum_1_cr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(611), ack => array_obj_ref_962_index_sum_1_req_1); -- 
    -- CP-element group 612 transition  input  output  no-bypass 
    -- predecessors 611 
    -- successors 613 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_index_sum_1_ack_1, ack => cp_elements(612)); -- 
    final_index_req_3390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(612), ack => array_obj_ref_962_offset_inst_req_0); -- 
    -- CP-element group 613 transition  input  output  no-bypass 
    -- predecessors 612 
    -- successors 614 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_offset_inst_ack_0, ack => cp_elements(613)); -- 
    sum_rename_req_3395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(613), ack => array_obj_ref_962_root_address_inst_req_0); -- 
    -- CP-element group 614 transition  input  no-bypass 
    -- predecessors 613 
    -- successors 601 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_962_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_962_root_address_inst_ack_0, ack => cp_elements(614)); -- 
    -- CP-element group 615 transition  output  bypass 
    -- predecessors 601 
    -- successors 616 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_963_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_963_complete/final_reg_req
      -- 
    cp_elements(615) <= cp_elements(601);
    final_reg_req_3400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(615), ack => addr_of_963_final_reg_req_0); -- 
    -- CP-element group 616 transition  input  no-bypass 
    -- predecessors 615 
    -- successors 602 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_963_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_963_complete/final_reg_ack
      -- 
    final_reg_ack_3401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_963_final_reg_ack_0, ack => cp_elements(616)); -- 
    -- CP-element group 617 transition  bypass 
    -- predecessors 367 
    -- successors 618 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_969_trigger_
      -- 
    cp_elements(617) <= cp_elements(367);
    -- CP-element group 618 join  fork  transition  no-bypass 
    -- predecessors 617 631 
    -- successors 619 632 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_969_active_
      -- 
    cpelement_group_618 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(617);
      predecessors(1) <= cp_elements(631);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(618)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(618),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 619 join  transition  output  bypass 
    -- predecessors 618 633 
    -- successors 1450 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_970_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_970_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_970_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_969_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1352_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1352_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1352_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_addr_resize/base_resize_req
      -- 
    cpelement_group_619 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(618);
      predecessors(1) <= cp_elements(633);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(619)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(619),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_6482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(619), ack => ptr_deref_1353_base_resize_req_0); -- 
    -- CP-element group 620 join  transition  output  bypass 
    -- predecessors 624 627 
    -- successors 628 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_620 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(624);
      predecessors(1) <= cp_elements(627);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(620)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(620),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(620), ack => array_obj_ref_968_index_sum_1_req_0); -- 
    -- CP-element group 621 transition  output  bypass 
    -- predecessors 367 
    -- successors 622 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_966_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_966_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_966_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_0/index_resize_req
      -- 
    cp_elements(621) <= cp_elements(367);
    index_resize_req_3419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(621), ack => array_obj_ref_968_index_0_resize_req_0); -- 
    -- CP-element group 622 transition  input  output  no-bypass 
    -- predecessors 621 
    -- successors 623 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_0/scale_rr
      -- 
    index_resize_ack_3420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_index_0_resize_ack_0, ack => cp_elements(622)); -- 
    scale_rr_3424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(622), ack => array_obj_ref_968_index_0_scale_req_0); -- 
    -- CP-element group 623 transition  input  output  no-bypass 
    -- predecessors 622 
    -- successors 624 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_0/scale_cr
      -- 
    scale_ra_3425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_index_0_scale_ack_0, ack => cp_elements(623)); -- 
    scale_cr_3426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(623), ack => array_obj_ref_968_index_0_scale_req_1); -- 
    -- CP-element group 624 transition  input  no-bypass 
    -- predecessors 623 
    -- successors 620 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_0/scale_ca
      -- 
    scale_ca_3427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_index_0_scale_ack_1, ack => cp_elements(624)); -- 
    -- CP-element group 625 transition  output  bypass 
    -- predecessors 417 
    -- successors 626 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_967_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_967_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_967_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_1/index_resize_req
      -- 
    cp_elements(625) <= cp_elements(417);
    index_resize_req_3436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(625), ack => array_obj_ref_968_index_1_resize_req_0); -- 
    -- CP-element group 626 transition  input  output  no-bypass 
    -- predecessors 625 
    -- successors 627 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_index_1_resize_ack_0, ack => cp_elements(626)); -- 
    scale_rename_req_3441_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(626), ack => array_obj_ref_968_index_1_rename_req_0); -- 
    -- CP-element group 627 transition  input  no-bypass 
    -- predecessors 626 
    -- successors 620 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3442_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_index_1_rename_ack_0, ack => cp_elements(627)); -- 
    -- CP-element group 628 transition  input  output  no-bypass 
    -- predecessors 620 
    -- successors 629 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3447_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_index_sum_1_ack_0, ack => cp_elements(628)); -- 
    partial_sum_1_cr_3448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(628), ack => array_obj_ref_968_index_sum_1_req_1); -- 
    -- CP-element group 629 transition  input  output  no-bypass 
    -- predecessors 628 
    -- successors 630 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_index_sum_1_ack_1, ack => cp_elements(629)); -- 
    final_index_req_3450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(629), ack => array_obj_ref_968_offset_inst_req_0); -- 
    -- CP-element group 630 transition  input  output  no-bypass 
    -- predecessors 629 
    -- successors 631 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_offset_inst_ack_0, ack => cp_elements(630)); -- 
    sum_rename_req_3455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(630), ack => array_obj_ref_968_root_address_inst_req_0); -- 
    -- CP-element group 631 transition  input  no-bypass 
    -- predecessors 630 
    -- successors 618 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_968_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_968_root_address_inst_ack_0, ack => cp_elements(631)); -- 
    -- CP-element group 632 transition  output  bypass 
    -- predecessors 618 
    -- successors 633 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_969_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_969_complete/final_reg_req
      -- 
    cp_elements(632) <= cp_elements(618);
    final_reg_req_3460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(632), ack => addr_of_969_final_reg_req_0); -- 
    -- CP-element group 633 transition  input  no-bypass 
    -- predecessors 632 
    -- successors 619 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_969_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_969_complete/final_reg_ack
      -- 
    final_reg_ack_3461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_969_final_reg_ack_0, ack => cp_elements(633)); -- 
    -- CP-element group 634 transition  bypass 
    -- predecessors 367 
    -- successors 635 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_975_trigger_
      -- 
    cp_elements(634) <= cp_elements(367);
    -- CP-element group 635 join  fork  transition  no-bypass 
    -- predecessors 634 648 
    -- successors 636 649 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_975_active_
      -- 
    cpelement_group_635 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(634);
      predecessors(1) <= cp_elements(648);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(635)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(635),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 636 join  transition  output  bypass 
    -- predecessors 635 650 
    -- successors 1440 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_976_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_976_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_976_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_975_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1348_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1348_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1348_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_addr_resize/base_resize_req
      -- 
    cpelement_group_636 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(635);
      predecessors(1) <= cp_elements(650);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(636)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(636),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_6430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => ptr_deref_1349_base_resize_req_0); -- 
    -- CP-element group 637 join  transition  output  bypass 
    -- predecessors 641 644 
    -- successors 645 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_637 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(641);
      predecessors(1) <= cp_elements(644);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(637)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(637),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3506_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(637), ack => array_obj_ref_974_index_sum_1_req_0); -- 
    -- CP-element group 638 transition  output  bypass 
    -- predecessors 367 
    -- successors 639 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_972_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_972_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_972_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_0/index_resize_req
      -- 
    cp_elements(638) <= cp_elements(367);
    index_resize_req_3479_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(638), ack => array_obj_ref_974_index_0_resize_req_0); -- 
    -- CP-element group 639 transition  input  output  no-bypass 
    -- predecessors 638 
    -- successors 640 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_0/scale_rr
      -- 
    index_resize_ack_3480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_index_0_resize_ack_0, ack => cp_elements(639)); -- 
    scale_rr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(639), ack => array_obj_ref_974_index_0_scale_req_0); -- 
    -- CP-element group 640 transition  input  output  no-bypass 
    -- predecessors 639 
    -- successors 641 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_0/scale_cr
      -- 
    scale_ra_3485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_index_0_scale_ack_0, ack => cp_elements(640)); -- 
    scale_cr_3486_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(640), ack => array_obj_ref_974_index_0_scale_req_1); -- 
    -- CP-element group 641 transition  input  no-bypass 
    -- predecessors 640 
    -- successors 637 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_0/scale_ca
      -- 
    scale_ca_3487_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_index_0_scale_ack_1, ack => cp_elements(641)); -- 
    -- CP-element group 642 transition  output  bypass 
    -- predecessors 492 
    -- successors 643 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_973_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_973_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_973_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_1/index_resize_req
      -- 
    cp_elements(642) <= cp_elements(492);
    index_resize_req_3496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(642), ack => array_obj_ref_974_index_1_resize_req_0); -- 
    -- CP-element group 643 transition  input  output  no-bypass 
    -- predecessors 642 
    -- successors 644 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_index_1_resize_ack_0, ack => cp_elements(643)); -- 
    scale_rename_req_3501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(643), ack => array_obj_ref_974_index_1_rename_req_0); -- 
    -- CP-element group 644 transition  input  no-bypass 
    -- predecessors 643 
    -- successors 637 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_index_1_rename_ack_0, ack => cp_elements(644)); -- 
    -- CP-element group 645 transition  input  output  no-bypass 
    -- predecessors 637 
    -- successors 646 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3507_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_index_sum_1_ack_0, ack => cp_elements(645)); -- 
    partial_sum_1_cr_3508_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(645), ack => array_obj_ref_974_index_sum_1_req_1); -- 
    -- CP-element group 646 transition  input  output  no-bypass 
    -- predecessors 645 
    -- successors 647 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3509_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_index_sum_1_ack_1, ack => cp_elements(646)); -- 
    final_index_req_3510_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(646), ack => array_obj_ref_974_offset_inst_req_0); -- 
    -- CP-element group 647 transition  input  output  no-bypass 
    -- predecessors 646 
    -- successors 648 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3511_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_offset_inst_ack_0, ack => cp_elements(647)); -- 
    sum_rename_req_3515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(647), ack => array_obj_ref_974_root_address_inst_req_0); -- 
    -- CP-element group 648 transition  input  no-bypass 
    -- predecessors 647 
    -- successors 635 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_974_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_974_root_address_inst_ack_0, ack => cp_elements(648)); -- 
    -- CP-element group 649 transition  output  bypass 
    -- predecessors 635 
    -- successors 650 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_975_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_975_complete/final_reg_req
      -- 
    cp_elements(649) <= cp_elements(635);
    final_reg_req_3520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(649), ack => addr_of_975_final_reg_req_0); -- 
    -- CP-element group 650 transition  input  no-bypass 
    -- predecessors 649 
    -- successors 636 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_975_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_975_complete/final_reg_ack
      -- 
    final_reg_ack_3521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_975_final_reg_ack_0, ack => cp_elements(650)); -- 
    -- CP-element group 651 transition  bypass 
    -- predecessors 367 
    -- successors 652 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_981_trigger_
      -- 
    cp_elements(651) <= cp_elements(367);
    -- CP-element group 652 join  fork  transition  no-bypass 
    -- predecessors 651 665 
    -- successors 653 666 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_981_active_
      -- 
    cpelement_group_652 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(651);
      predecessors(1) <= cp_elements(665);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(652)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(652),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 653 join  transition  output  bypass 
    -- predecessors 652 667 
    -- successors 990 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_982_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_982_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_982_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_981_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1112_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1112_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1112_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_addr_resize/base_resize_req
      -- 
    cpelement_group_653 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(652);
      predecessors(1) <= cp_elements(667);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(653)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(653),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(653), ack => ptr_deref_1113_base_resize_req_0); -- 
    -- CP-element group 654 join  transition  output  bypass 
    -- predecessors 658 661 
    -- successors 662 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_654 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(658);
      predecessors(1) <= cp_elements(661);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(654)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(654),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => array_obj_ref_980_index_sum_1_req_0); -- 
    -- CP-element group 655 transition  output  bypass 
    -- predecessors 367 
    -- successors 656 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_978_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_978_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_978_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_0/index_resize_req
      -- 
    cp_elements(655) <= cp_elements(367);
    index_resize_req_3539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(655), ack => array_obj_ref_980_index_0_resize_req_0); -- 
    -- CP-element group 656 transition  input  output  no-bypass 
    -- predecessors 655 
    -- successors 657 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_0/scale_rr
      -- 
    index_resize_ack_3540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_index_0_resize_ack_0, ack => cp_elements(656)); -- 
    scale_rr_3544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(656), ack => array_obj_ref_980_index_0_scale_req_0); -- 
    -- CP-element group 657 transition  input  output  no-bypass 
    -- predecessors 656 
    -- successors 658 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_0/scale_cr
      -- 
    scale_ra_3545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_index_0_scale_ack_0, ack => cp_elements(657)); -- 
    scale_cr_3546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(657), ack => array_obj_ref_980_index_0_scale_req_1); -- 
    -- CP-element group 658 transition  input  no-bypass 
    -- predecessors 657 
    -- successors 654 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_0/scale_ca
      -- 
    scale_ca_3547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_index_0_scale_ack_1, ack => cp_elements(658)); -- 
    -- CP-element group 659 transition  output  bypass 
    -- predecessors 492 
    -- successors 660 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_979_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_979_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_979_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_1/index_resize_req
      -- 
    cp_elements(659) <= cp_elements(492);
    index_resize_req_3556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(659), ack => array_obj_ref_980_index_1_resize_req_0); -- 
    -- CP-element group 660 transition  input  output  no-bypass 
    -- predecessors 659 
    -- successors 661 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_index_1_resize_ack_0, ack => cp_elements(660)); -- 
    scale_rename_req_3561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(660), ack => array_obj_ref_980_index_1_rename_req_0); -- 
    -- CP-element group 661 transition  input  no-bypass 
    -- predecessors 660 
    -- successors 654 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_index_1_rename_ack_0, ack => cp_elements(661)); -- 
    -- CP-element group 662 transition  input  output  no-bypass 
    -- predecessors 654 
    -- successors 663 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_index_sum_1_ack_0, ack => cp_elements(662)); -- 
    partial_sum_1_cr_3568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(662), ack => array_obj_ref_980_index_sum_1_req_1); -- 
    -- CP-element group 663 transition  input  output  no-bypass 
    -- predecessors 662 
    -- successors 664 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_index_sum_1_ack_1, ack => cp_elements(663)); -- 
    final_index_req_3570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(663), ack => array_obj_ref_980_offset_inst_req_0); -- 
    -- CP-element group 664 transition  input  output  no-bypass 
    -- predecessors 663 
    -- successors 665 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_offset_inst_ack_0, ack => cp_elements(664)); -- 
    sum_rename_req_3575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(664), ack => array_obj_ref_980_root_address_inst_req_0); -- 
    -- CP-element group 665 transition  input  no-bypass 
    -- predecessors 664 
    -- successors 652 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_980_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_980_root_address_inst_ack_0, ack => cp_elements(665)); -- 
    -- CP-element group 666 transition  output  bypass 
    -- predecessors 652 
    -- successors 667 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_981_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_981_complete/final_reg_req
      -- 
    cp_elements(666) <= cp_elements(652);
    final_reg_req_3580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(666), ack => addr_of_981_final_reg_req_0); -- 
    -- CP-element group 667 transition  input  no-bypass 
    -- predecessors 666 
    -- successors 653 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_981_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_981_complete/final_reg_ack
      -- 
    final_reg_ack_3581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_981_final_reg_ack_0, ack => cp_elements(667)); -- 
    -- CP-element group 668 join  fork  transition  no-bypass 
    -- predecessors 670 672 
    -- successors 669 673 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_active_
      -- 
    cpelement_group_668 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(670);
      predecessors(1) <= cp_elements(672);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(668)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(668),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 669 join  fork  transition  bypass 
    -- predecessors 668 674 
    -- successors 677 701 725 751 819 887 955 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_988_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_988_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_988_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_completed_
      -- 
    cpelement_group_669 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(668);
      predecessors(1) <= cp_elements(674);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(669)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(669),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 670 fork  transition  bypass 
    -- predecessors 367 
    -- successors 668 671 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_984_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_984_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_984_completed_
      -- 
    cp_elements(670) <= cp_elements(367);
    -- CP-element group 671 transition  output  bypass 
    -- predecessors 670 
    -- successors 672 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Sample/rr
      -- 
    cp_elements(671) <= cp_elements(670);
    rr_3594_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(671), ack => binary_987_inst_req_0); -- 
    -- CP-element group 672 transition  input  no-bypass 
    -- predecessors 671 
    -- successors 668 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Sample/ra
      -- 
    ra_3595_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_987_inst_ack_0, ack => cp_elements(672)); -- 
    -- CP-element group 673 transition  output  bypass 
    -- predecessors 668 
    -- successors 674 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Update/cr
      -- 
    cp_elements(673) <= cp_elements(668);
    cr_3599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(673), ack => binary_987_inst_req_1); -- 
    -- CP-element group 674 transition  input  no-bypass 
    -- predecessors 673 
    -- successors 669 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_987_complete_Update/ca
      -- 
    ca_3600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_987_inst_ack_1, ack => cp_elements(674)); -- 
    -- CP-element group 675 join  fork  transition  no-bypass 
    -- predecessors 677 679 
    -- successors 676 680 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_active_
      -- 
    cpelement_group_675 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(677);
      predecessors(1) <= cp_elements(679);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(675)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(675),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 676 join  fork  transition  no-bypass 
    -- predecessors 675 681 
    -- successors 686 768 836 904 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_994_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_994_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_994_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_completed_
      -- 
    cpelement_group_676 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(675);
      predecessors(1) <= cp_elements(681);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(676)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(676),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 677 fork  transition  bypass 
    -- predecessors 669 
    -- successors 675 678 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_990_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_990_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_990_completed_
      -- 
    cp_elements(677) <= cp_elements(669);
    -- CP-element group 678 transition  output  bypass 
    -- predecessors 677 
    -- successors 679 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Sample/rr
      -- 
    cp_elements(678) <= cp_elements(677);
    rr_3613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(678), ack => binary_993_inst_req_0); -- 
    -- CP-element group 679 transition  input  no-bypass 
    -- predecessors 678 
    -- successors 675 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Sample/ra
      -- 
    ra_3614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_993_inst_ack_0, ack => cp_elements(679)); -- 
    -- CP-element group 680 transition  output  bypass 
    -- predecessors 675 
    -- successors 681 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Update/cr
      -- 
    cp_elements(680) <= cp_elements(675);
    cr_3618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(680), ack => binary_993_inst_req_1); -- 
    -- CP-element group 681 transition  input  no-bypass 
    -- predecessors 680 
    -- successors 676 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_993_complete_Update/ca
      -- 
    ca_3619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_993_inst_ack_1, ack => cp_elements(681)); -- 
    -- CP-element group 682 transition  bypass 
    -- predecessors 367 
    -- successors 683 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_999_trigger_
      -- 
    cp_elements(682) <= cp_elements(367);
    -- CP-element group 683 join  fork  transition  no-bypass 
    -- predecessors 682 696 
    -- successors 684 697 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_999_active_
      -- 
    cpelement_group_683 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(682);
      predecessors(1) <= cp_elements(696);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(683)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(683),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 684 join  transition  output  bypass 
    -- predecessors 683 698 
    -- successors 1040 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1000_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1000_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1000_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_999_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1132_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1132_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1132_completed_
      -- 
    cpelement_group_684 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(683);
      predecessors(1) <= cp_elements(698);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(684)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(684),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(684), ack => ptr_deref_1133_base_resize_req_0); -- 
    -- CP-element group 685 join  transition  output  bypass 
    -- predecessors 689 692 
    -- successors 693 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_685 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(689);
      predecessors(1) <= cp_elements(692);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(685)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(685),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(685), ack => array_obj_ref_998_index_sum_1_req_0); -- 
    -- CP-element group 686 transition  output  bypass 
    -- predecessors 676 
    -- successors 687 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_996_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_996_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_996_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_0/index_resize_req
      -- 
    cp_elements(686) <= cp_elements(676);
    index_resize_req_3637_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(686), ack => array_obj_ref_998_index_0_resize_req_0); -- 
    -- CP-element group 687 transition  input  output  no-bypass 
    -- predecessors 686 
    -- successors 688 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_0/scale_rr
      -- 
    index_resize_ack_3638_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_0_resize_ack_0, ack => cp_elements(687)); -- 
    scale_rr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(687), ack => array_obj_ref_998_index_0_scale_req_0); -- 
    -- CP-element group 688 transition  input  output  no-bypass 
    -- predecessors 687 
    -- successors 689 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_0/scale_cr
      -- 
    scale_ra_3643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_0_scale_ack_0, ack => cp_elements(688)); -- 
    scale_cr_3644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(688), ack => array_obj_ref_998_index_0_scale_req_1); -- 
    -- CP-element group 689 transition  input  no-bypass 
    -- predecessors 688 
    -- successors 685 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_0/scale_ca
      -- 
    scale_ca_3645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_0_scale_ack_1, ack => cp_elements(689)); -- 
    -- CP-element group 690 transition  output  bypass 
    -- predecessors 367 
    -- successors 691 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_997_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_997_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_997_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_1/index_resize_req
      -- 
    cp_elements(690) <= cp_elements(367);
    index_resize_req_3654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => array_obj_ref_998_index_1_resize_req_0); -- 
    -- CP-element group 691 transition  input  output  no-bypass 
    -- predecessors 690 
    -- successors 692 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_1_resize_ack_0, ack => cp_elements(691)); -- 
    scale_rename_req_3659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(691), ack => array_obj_ref_998_index_1_rename_req_0); -- 
    -- CP-element group 692 transition  input  no-bypass 
    -- predecessors 691 
    -- successors 685 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_1_rename_ack_0, ack => cp_elements(692)); -- 
    -- CP-element group 693 transition  input  output  no-bypass 
    -- predecessors 685 
    -- successors 694 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_sum_1_ack_0, ack => cp_elements(693)); -- 
    partial_sum_1_cr_3666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(693), ack => array_obj_ref_998_index_sum_1_req_1); -- 
    -- CP-element group 694 transition  input  output  no-bypass 
    -- predecessors 693 
    -- successors 695 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_index_sum_1_ack_1, ack => cp_elements(694)); -- 
    final_index_req_3668_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => array_obj_ref_998_offset_inst_req_0); -- 
    -- CP-element group 695 transition  input  output  no-bypass 
    -- predecessors 694 
    -- successors 696 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3669_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_offset_inst_ack_0, ack => cp_elements(695)); -- 
    sum_rename_req_3673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(695), ack => array_obj_ref_998_root_address_inst_req_0); -- 
    -- CP-element group 696 transition  input  no-bypass 
    -- predecessors 695 
    -- successors 683 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_998_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3674_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_998_root_address_inst_ack_0, ack => cp_elements(696)); -- 
    -- CP-element group 697 transition  output  bypass 
    -- predecessors 683 
    -- successors 698 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_999_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_999_complete/final_reg_req
      -- 
    cp_elements(697) <= cp_elements(683);
    final_reg_req_3678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(697), ack => addr_of_999_final_reg_req_0); -- 
    -- CP-element group 698 transition  input  no-bypass 
    -- predecessors 697 
    -- successors 684 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_999_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_999_complete/final_reg_ack
      -- 
    final_reg_ack_3679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_999_final_reg_ack_0, ack => cp_elements(698)); -- 
    -- CP-element group 699 join  fork  transition  no-bypass 
    -- predecessors 701 703 
    -- successors 700 704 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_active_
      -- 
    cpelement_group_699 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(701);
      predecessors(1) <= cp_elements(703);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(699)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(699),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 700 join  fork  transition  no-bypass 
    -- predecessors 699 705 
    -- successors 710 785 853 921 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1006_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1006_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1006_completed_
      -- 
    cpelement_group_700 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(699);
      predecessors(1) <= cp_elements(705);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(700)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(700),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 701 fork  transition  bypass 
    -- predecessors 669 
    -- successors 699 702 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1002_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1002_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1002_completed_
      -- 
    cp_elements(701) <= cp_elements(669);
    -- CP-element group 702 transition  output  bypass 
    -- predecessors 701 
    -- successors 703 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Sample/rr
      -- 
    cp_elements(702) <= cp_elements(701);
    rr_3692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(702), ack => binary_1005_inst_req_0); -- 
    -- CP-element group 703 transition  input  no-bypass 
    -- predecessors 702 
    -- successors 699 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Sample/ra
      -- 
    ra_3693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1005_inst_ack_0, ack => cp_elements(703)); -- 
    -- CP-element group 704 transition  output  bypass 
    -- predecessors 699 
    -- successors 705 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Update/cr
      -- 
    cp_elements(704) <= cp_elements(699);
    cr_3697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(704), ack => binary_1005_inst_req_1); -- 
    -- CP-element group 705 transition  input  no-bypass 
    -- predecessors 704 
    -- successors 700 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1005_complete_Update/ca
      -- 
    ca_3698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1005_inst_ack_1, ack => cp_elements(705)); -- 
    -- CP-element group 706 transition  bypass 
    -- predecessors 367 
    -- successors 707 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1011_trigger_
      -- 
    cp_elements(706) <= cp_elements(367);
    -- CP-element group 707 join  fork  transition  no-bypass 
    -- predecessors 706 720 
    -- successors 708 721 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1011_active_
      -- 
    cpelement_group_707 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(706);
      predecessors(1) <= cp_elements(720);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(707)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(707),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 708 join  transition  output  bypass 
    -- predecessors 707 722 
    -- successors 1020 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1012_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1012_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1012_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1011_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1124_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1124_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1124_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_addr_resize/base_resize_req
      -- 
    cpelement_group_708 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(707);
      predecessors(1) <= cp_elements(722);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(708)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(708),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(708), ack => ptr_deref_1125_base_resize_req_0); -- 
    -- CP-element group 709 join  transition  output  bypass 
    -- predecessors 713 716 
    -- successors 717 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_709 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(713);
      predecessors(1) <= cp_elements(716);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(709)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(709),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(709), ack => array_obj_ref_1010_index_sum_1_req_0); -- 
    -- CP-element group 710 transition  output  bypass 
    -- predecessors 700 
    -- successors 711 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1008_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1008_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1008_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_0/index_resize_req
      -- 
    cp_elements(710) <= cp_elements(700);
    index_resize_req_3716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(710), ack => array_obj_ref_1010_index_0_resize_req_0); -- 
    -- CP-element group 711 transition  input  output  no-bypass 
    -- predecessors 710 
    -- successors 712 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_0/scale_rr
      -- 
    index_resize_ack_3717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_index_0_resize_ack_0, ack => cp_elements(711)); -- 
    scale_rr_3721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => array_obj_ref_1010_index_0_scale_req_0); -- 
    -- CP-element group 712 transition  input  output  no-bypass 
    -- predecessors 711 
    -- successors 713 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_0/scale_cr
      -- 
    scale_ra_3722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_index_0_scale_ack_0, ack => cp_elements(712)); -- 
    scale_cr_3723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(712), ack => array_obj_ref_1010_index_0_scale_req_1); -- 
    -- CP-element group 713 transition  input  no-bypass 
    -- predecessors 712 
    -- successors 709 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_0/scale_ca
      -- 
    scale_ca_3724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_index_0_scale_ack_1, ack => cp_elements(713)); -- 
    -- CP-element group 714 transition  output  bypass 
    -- predecessors 367 
    -- successors 715 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1009_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1009_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1009_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_1/index_resize_req
      -- 
    cp_elements(714) <= cp_elements(367);
    index_resize_req_3733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(714), ack => array_obj_ref_1010_index_1_resize_req_0); -- 
    -- CP-element group 715 transition  input  output  no-bypass 
    -- predecessors 714 
    -- successors 716 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_index_1_resize_ack_0, ack => cp_elements(715)); -- 
    scale_rename_req_3738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(715), ack => array_obj_ref_1010_index_1_rename_req_0); -- 
    -- CP-element group 716 transition  input  no-bypass 
    -- predecessors 715 
    -- successors 709 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3739_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_index_1_rename_ack_0, ack => cp_elements(716)); -- 
    -- CP-element group 717 transition  input  output  no-bypass 
    -- predecessors 709 
    -- successors 718 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_index_sum_1_ack_0, ack => cp_elements(717)); -- 
    partial_sum_1_cr_3745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(717), ack => array_obj_ref_1010_index_sum_1_req_1); -- 
    -- CP-element group 718 transition  input  output  no-bypass 
    -- predecessors 717 
    -- successors 719 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_index_sum_1_ack_1, ack => cp_elements(718)); -- 
    final_index_req_3747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(718), ack => array_obj_ref_1010_offset_inst_req_0); -- 
    -- CP-element group 719 transition  input  output  no-bypass 
    -- predecessors 718 
    -- successors 720 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_offset_inst_ack_0, ack => cp_elements(719)); -- 
    sum_rename_req_3752_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(719), ack => array_obj_ref_1010_root_address_inst_req_0); -- 
    -- CP-element group 720 transition  input  no-bypass 
    -- predecessors 719 
    -- successors 707 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1010_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3753_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1010_root_address_inst_ack_0, ack => cp_elements(720)); -- 
    -- CP-element group 721 transition  output  bypass 
    -- predecessors 707 
    -- successors 722 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1011_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1011_complete/final_reg_req
      -- 
    cp_elements(721) <= cp_elements(707);
    final_reg_req_3757_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(721), ack => addr_of_1011_final_reg_req_0); -- 
    -- CP-element group 722 transition  input  no-bypass 
    -- predecessors 721 
    -- successors 708 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1011_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1011_complete/final_reg_ack
      -- 
    final_reg_ack_3758_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1011_final_reg_ack_0, ack => cp_elements(722)); -- 
    -- CP-element group 723 join  fork  transition  no-bypass 
    -- predecessors 725 727 
    -- successors 724 728 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_active_
      -- 
    cpelement_group_723 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(725);
      predecessors(1) <= cp_elements(727);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(723)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(723),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 724 join  fork  transition  no-bypass 
    -- predecessors 723 729 
    -- successors 734 802 870 938 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1018_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1018_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1018_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_completed_
      -- 
    cpelement_group_724 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(723);
      predecessors(1) <= cp_elements(729);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(724)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(724),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 725 fork  transition  bypass 
    -- predecessors 669 
    -- successors 723 726 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1014_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1014_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1014_completed_
      -- 
    cp_elements(725) <= cp_elements(669);
    -- CP-element group 726 transition  output  bypass 
    -- predecessors 725 
    -- successors 727 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Sample/rr
      -- 
    cp_elements(726) <= cp_elements(725);
    rr_3771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(726), ack => binary_1017_inst_req_0); -- 
    -- CP-element group 727 transition  input  no-bypass 
    -- predecessors 726 
    -- successors 723 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Sample/ra
      -- 
    ra_3772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1017_inst_ack_0, ack => cp_elements(727)); -- 
    -- CP-element group 728 transition  output  bypass 
    -- predecessors 723 
    -- successors 729 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Update/cr
      -- 
    cp_elements(728) <= cp_elements(723);
    cr_3776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(728), ack => binary_1017_inst_req_1); -- 
    -- CP-element group 729 transition  input  no-bypass 
    -- predecessors 728 
    -- successors 724 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1017_complete_Update/ca
      -- 
    ca_3777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1017_inst_ack_1, ack => cp_elements(729)); -- 
    -- CP-element group 730 transition  bypass 
    -- predecessors 367 
    -- successors 731 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1023_trigger_
      -- 
    cp_elements(730) <= cp_elements(367);
    -- CP-element group 731 join  fork  transition  no-bypass 
    -- predecessors 730 744 
    -- successors 732 745 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1023_active_
      -- 
    cpelement_group_731 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(730);
      predecessors(1) <= cp_elements(744);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(731)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(731),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 732 join  transition  output  bypass 
    -- predecessors 731 746 
    -- successors 1000 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1024_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1024_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1024_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1023_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1116_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1116_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1116_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_addr_resize/base_resize_req
      -- 
    cpelement_group_732 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(731);
      predecessors(1) <= cp_elements(746);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(732)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(732),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(732), ack => ptr_deref_1117_base_resize_req_0); -- 
    -- CP-element group 733 join  transition  output  bypass 
    -- predecessors 737 740 
    -- successors 741 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_733 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(737);
      predecessors(1) <= cp_elements(740);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(733)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(733),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(733), ack => array_obj_ref_1022_index_sum_1_req_0); -- 
    -- CP-element group 734 transition  output  bypass 
    -- predecessors 724 
    -- successors 735 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1020_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1020_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1020_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_0/index_resize_req
      -- 
    cp_elements(734) <= cp_elements(724);
    index_resize_req_3795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(734), ack => array_obj_ref_1022_index_0_resize_req_0); -- 
    -- CP-element group 735 transition  input  output  no-bypass 
    -- predecessors 734 
    -- successors 736 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_0/scale_rr
      -- 
    index_resize_ack_3796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_index_0_resize_ack_0, ack => cp_elements(735)); -- 
    scale_rr_3800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => array_obj_ref_1022_index_0_scale_req_0); -- 
    -- CP-element group 736 transition  input  output  no-bypass 
    -- predecessors 735 
    -- successors 737 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_0/scale_cr
      -- 
    scale_ra_3801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_index_0_scale_ack_0, ack => cp_elements(736)); -- 
    scale_cr_3802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(736), ack => array_obj_ref_1022_index_0_scale_req_1); -- 
    -- CP-element group 737 transition  input  no-bypass 
    -- predecessors 736 
    -- successors 733 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_0/scale_ca
      -- 
    scale_ca_3803_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_index_0_scale_ack_1, ack => cp_elements(737)); -- 
    -- CP-element group 738 transition  output  bypass 
    -- predecessors 367 
    -- successors 739 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1021_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1021_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1021_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_1/index_resize_req
      -- 
    cp_elements(738) <= cp_elements(367);
    index_resize_req_3812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(738), ack => array_obj_ref_1022_index_1_resize_req_0); -- 
    -- CP-element group 739 transition  input  output  no-bypass 
    -- predecessors 738 
    -- successors 740 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_index_1_resize_ack_0, ack => cp_elements(739)); -- 
    scale_rename_req_3817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(739), ack => array_obj_ref_1022_index_1_rename_req_0); -- 
    -- CP-element group 740 transition  input  no-bypass 
    -- predecessors 739 
    -- successors 733 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_index_1_rename_ack_0, ack => cp_elements(740)); -- 
    -- CP-element group 741 transition  input  output  no-bypass 
    -- predecessors 733 
    -- successors 742 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_index_sum_1_ack_0, ack => cp_elements(741)); -- 
    partial_sum_1_cr_3824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(741), ack => array_obj_ref_1022_index_sum_1_req_1); -- 
    -- CP-element group 742 transition  input  output  no-bypass 
    -- predecessors 741 
    -- successors 743 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_index_sum_1_ack_1, ack => cp_elements(742)); -- 
    final_index_req_3826_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(742), ack => array_obj_ref_1022_offset_inst_req_0); -- 
    -- CP-element group 743 transition  input  output  no-bypass 
    -- predecessors 742 
    -- successors 744 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_offset_inst_ack_0, ack => cp_elements(743)); -- 
    sum_rename_req_3831_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(743), ack => array_obj_ref_1022_root_address_inst_req_0); -- 
    -- CP-element group 744 transition  input  no-bypass 
    -- predecessors 743 
    -- successors 731 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1022_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3832_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1022_root_address_inst_ack_0, ack => cp_elements(744)); -- 
    -- CP-element group 745 transition  output  bypass 
    -- predecessors 731 
    -- successors 746 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1023_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1023_complete/final_reg_req
      -- 
    cp_elements(745) <= cp_elements(731);
    final_reg_req_3836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(745), ack => addr_of_1023_final_reg_req_0); -- 
    -- CP-element group 746 transition  input  no-bypass 
    -- predecessors 745 
    -- successors 732 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1023_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1023_complete/final_reg_ack
      -- 
    final_reg_ack_3837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1023_final_reg_ack_0, ack => cp_elements(746)); -- 
    -- CP-element group 747 transition  bypass 
    -- predecessors 367 
    -- successors 748 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1029_trigger_
      -- 
    cp_elements(747) <= cp_elements(367);
    -- CP-element group 748 join  fork  transition  no-bypass 
    -- predecessors 747 761 
    -- successors 749 762 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1029_active_
      -- 
    cpelement_group_748 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(747);
      predecessors(1) <= cp_elements(761);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(748)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(748),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 749 join  transition  output  bypass 
    -- predecessors 748 763 
    -- successors 980 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1030_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1030_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1030_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1029_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1108_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1108_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1108_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_addr_resize/base_resize_req
      -- 
    cpelement_group_749 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(748);
      predecessors(1) <= cp_elements(763);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(749)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(749),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_4686_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(749), ack => ptr_deref_1109_base_resize_req_0); -- 
    -- CP-element group 750 join  transition  output  bypass 
    -- predecessors 754 757 
    -- successors 758 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_750 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(754);
      predecessors(1) <= cp_elements(757);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(750)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(750),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(750), ack => array_obj_ref_1028_index_sum_1_req_0); -- 
    -- CP-element group 751 transition  output  bypass 
    -- predecessors 669 
    -- successors 752 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1026_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1026_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1026_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_0/index_resize_req
      -- 
    cp_elements(751) <= cp_elements(669);
    index_resize_req_3855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(751), ack => array_obj_ref_1028_index_0_resize_req_0); -- 
    -- CP-element group 752 transition  input  output  no-bypass 
    -- predecessors 751 
    -- successors 753 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_0/scale_rr
      -- 
    index_resize_ack_3856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_0_resize_ack_0, ack => cp_elements(752)); -- 
    scale_rr_3860_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(752), ack => array_obj_ref_1028_index_0_scale_req_0); -- 
    -- CP-element group 753 transition  input  output  no-bypass 
    -- predecessors 752 
    -- successors 754 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_0/scale_cr
      -- 
    scale_ra_3861_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_0_scale_ack_0, ack => cp_elements(753)); -- 
    scale_cr_3862_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(753), ack => array_obj_ref_1028_index_0_scale_req_1); -- 
    -- CP-element group 754 transition  input  no-bypass 
    -- predecessors 753 
    -- successors 750 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_0/scale_ca
      -- 
    scale_ca_3863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_0_scale_ack_1, ack => cp_elements(754)); -- 
    -- CP-element group 755 transition  output  bypass 
    -- predecessors 367 
    -- successors 756 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1027_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1027_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1027_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_1/index_resize_req
      -- 
    cp_elements(755) <= cp_elements(367);
    index_resize_req_3872_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(755), ack => array_obj_ref_1028_index_1_resize_req_0); -- 
    -- CP-element group 756 transition  input  output  no-bypass 
    -- predecessors 755 
    -- successors 757 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3873_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_1_resize_ack_0, ack => cp_elements(756)); -- 
    scale_rename_req_3877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => array_obj_ref_1028_index_1_rename_req_0); -- 
    -- CP-element group 757 transition  input  no-bypass 
    -- predecessors 756 
    -- successors 750 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_1_rename_ack_0, ack => cp_elements(757)); -- 
    -- CP-element group 758 transition  input  output  no-bypass 
    -- predecessors 750 
    -- successors 759 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3883_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_sum_1_ack_0, ack => cp_elements(758)); -- 
    partial_sum_1_cr_3884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(758), ack => array_obj_ref_1028_index_sum_1_req_1); -- 
    -- CP-element group 759 transition  input  output  no-bypass 
    -- predecessors 758 
    -- successors 760 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_index_sum_1_ack_1, ack => cp_elements(759)); -- 
    final_index_req_3886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(759), ack => array_obj_ref_1028_offset_inst_req_0); -- 
    -- CP-element group 760 transition  input  output  no-bypass 
    -- predecessors 759 
    -- successors 761 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_offset_inst_ack_0, ack => cp_elements(760)); -- 
    sum_rename_req_3891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(760), ack => array_obj_ref_1028_root_address_inst_req_0); -- 
    -- CP-element group 761 transition  input  no-bypass 
    -- predecessors 760 
    -- successors 748 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1028_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1028_root_address_inst_ack_0, ack => cp_elements(761)); -- 
    -- CP-element group 762 transition  output  bypass 
    -- predecessors 748 
    -- successors 763 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1029_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1029_complete/final_reg_req
      -- 
    cp_elements(762) <= cp_elements(748);
    final_reg_req_3896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(762), ack => addr_of_1029_final_reg_req_0); -- 
    -- CP-element group 763 transition  input  no-bypass 
    -- predecessors 762 
    -- successors 749 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1029_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1029_complete/final_reg_ack
      -- 
    final_reg_ack_3897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1029_final_reg_ack_0, ack => cp_elements(763)); -- 
    -- CP-element group 764 transition  bypass 
    -- predecessors 367 
    -- successors 765 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1035_trigger_
      -- 
    cp_elements(764) <= cp_elements(367);
    -- CP-element group 765 join  fork  transition  no-bypass 
    -- predecessors 764 778 
    -- successors 766 779 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1035_active_
      -- 
    cpelement_group_765 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(764);
      predecessors(1) <= cp_elements(778);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(765)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(765),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 766 join  transition  output  bypass 
    -- predecessors 765 780 
    -- successors 1145 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1036_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1036_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1036_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1035_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1188_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1188_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1188_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_addr_resize/base_resize_req
      -- 
    cpelement_group_766 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(765);
      predecessors(1) <= cp_elements(780);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(766)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(766),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(766), ack => ptr_deref_1189_base_resize_req_0); -- 
    -- CP-element group 767 join  transition  output  bypass 
    -- predecessors 771 774 
    -- successors 775 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_767 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(771);
      predecessors(1) <= cp_elements(774);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(767)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(767),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_3942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(767), ack => array_obj_ref_1034_index_sum_1_req_0); -- 
    -- CP-element group 768 transition  output  bypass 
    -- predecessors 676 
    -- successors 769 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1032_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1032_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1032_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_0/index_resize_req
      -- 
    cp_elements(768) <= cp_elements(676);
    index_resize_req_3915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(768), ack => array_obj_ref_1034_index_0_resize_req_0); -- 
    -- CP-element group 769 transition  input  output  no-bypass 
    -- predecessors 768 
    -- successors 770 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_0/scale_rr
      -- 
    index_resize_ack_3916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_0_resize_ack_0, ack => cp_elements(769)); -- 
    scale_rr_3920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(769), ack => array_obj_ref_1034_index_0_scale_req_0); -- 
    -- CP-element group 770 transition  input  output  no-bypass 
    -- predecessors 769 
    -- successors 771 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_0/scale_cr
      -- 
    scale_ra_3921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_0_scale_ack_0, ack => cp_elements(770)); -- 
    scale_cr_3922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(770), ack => array_obj_ref_1034_index_0_scale_req_1); -- 
    -- CP-element group 771 transition  input  no-bypass 
    -- predecessors 770 
    -- successors 767 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_0/scale_ca
      -- 
    scale_ca_3923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_0_scale_ack_1, ack => cp_elements(771)); -- 
    -- CP-element group 772 transition  output  bypass 
    -- predecessors 367 
    -- successors 773 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1033_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1033_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1033_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_1/index_resize_req
      -- 
    cp_elements(772) <= cp_elements(367);
    index_resize_req_3932_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(772), ack => array_obj_ref_1034_index_1_resize_req_0); -- 
    -- CP-element group 773 transition  input  output  no-bypass 
    -- predecessors 772 
    -- successors 774 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3933_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_1_resize_ack_0, ack => cp_elements(773)); -- 
    scale_rename_req_3937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(773), ack => array_obj_ref_1034_index_1_rename_req_0); -- 
    -- CP-element group 774 transition  input  no-bypass 
    -- predecessors 773 
    -- successors 767 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_1_rename_ack_0, ack => cp_elements(774)); -- 
    -- CP-element group 775 transition  input  output  no-bypass 
    -- predecessors 767 
    -- successors 776 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_3943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_sum_1_ack_0, ack => cp_elements(775)); -- 
    partial_sum_1_cr_3944_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(775), ack => array_obj_ref_1034_index_sum_1_req_1); -- 
    -- CP-element group 776 transition  input  output  no-bypass 
    -- predecessors 775 
    -- successors 777 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/final_index_req
      -- 
    partial_sum_1_ca_3945_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_index_sum_1_ack_1, ack => cp_elements(776)); -- 
    final_index_req_3946_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(776), ack => array_obj_ref_1034_offset_inst_req_0); -- 
    -- CP-element group 777 transition  input  output  no-bypass 
    -- predecessors 776 
    -- successors 778 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3947_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_offset_inst_ack_0, ack => cp_elements(777)); -- 
    sum_rename_req_3951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(777), ack => array_obj_ref_1034_root_address_inst_req_0); -- 
    -- CP-element group 778 transition  input  no-bypass 
    -- predecessors 777 
    -- successors 765 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1034_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1034_root_address_inst_ack_0, ack => cp_elements(778)); -- 
    -- CP-element group 779 transition  output  bypass 
    -- predecessors 765 
    -- successors 780 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1035_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1035_complete/final_reg_req
      -- 
    cp_elements(779) <= cp_elements(765);
    final_reg_req_3956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(779), ack => addr_of_1035_final_reg_req_0); -- 
    -- CP-element group 780 transition  input  no-bypass 
    -- predecessors 779 
    -- successors 766 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1035_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1035_complete/final_reg_ack
      -- 
    final_reg_ack_3957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1035_final_reg_ack_0, ack => cp_elements(780)); -- 
    -- CP-element group 781 transition  bypass 
    -- predecessors 367 
    -- successors 782 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1041_trigger_
      -- 
    cp_elements(781) <= cp_elements(367);
    -- CP-element group 782 join  fork  transition  no-bypass 
    -- predecessors 781 795 
    -- successors 783 796 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1041_active_
      -- 
    cpelement_group_782 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(781);
      predecessors(1) <= cp_elements(795);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(782)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(782),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 783 join  transition  output  bypass 
    -- predecessors 782 797 
    -- successors 1135 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1041_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1042_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1042_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1042_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1184_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1184_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1184_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_addr_resize/base_resize_req
      -- 
    cpelement_group_783 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(782);
      predecessors(1) <= cp_elements(797);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(783)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(783),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5330_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => ptr_deref_1185_base_resize_req_0); -- 
    -- CP-element group 784 join  transition  output  bypass 
    -- predecessors 788 791 
    -- successors 792 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_784 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(788);
      predecessors(1) <= cp_elements(791);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(784)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(784),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4002_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => array_obj_ref_1040_index_sum_1_req_0); -- 
    -- CP-element group 785 transition  output  bypass 
    -- predecessors 700 
    -- successors 786 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1038_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1038_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1038_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_0/index_resize_req
      -- 
    cp_elements(785) <= cp_elements(700);
    index_resize_req_3975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => array_obj_ref_1040_index_0_resize_req_0); -- 
    -- CP-element group 786 transition  input  output  no-bypass 
    -- predecessors 785 
    -- successors 787 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_0/scale_rr
      -- 
    index_resize_ack_3976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_0_resize_ack_0, ack => cp_elements(786)); -- 
    scale_rr_3980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(786), ack => array_obj_ref_1040_index_0_scale_req_0); -- 
    -- CP-element group 787 transition  input  output  no-bypass 
    -- predecessors 786 
    -- successors 788 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_0/scale_cr
      -- 
    scale_ra_3981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_0_scale_ack_0, ack => cp_elements(787)); -- 
    scale_cr_3982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(787), ack => array_obj_ref_1040_index_0_scale_req_1); -- 
    -- CP-element group 788 transition  input  no-bypass 
    -- predecessors 787 
    -- successors 784 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_0/scale_ca
      -- 
    scale_ca_3983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_0_scale_ack_1, ack => cp_elements(788)); -- 
    -- CP-element group 789 transition  output  bypass 
    -- predecessors 367 
    -- successors 790 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1039_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1039_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1039_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_1/index_resize_req
      -- 
    cp_elements(789) <= cp_elements(367);
    index_resize_req_3992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(789), ack => array_obj_ref_1040_index_1_resize_req_0); -- 
    -- CP-element group 790 transition  input  output  no-bypass 
    -- predecessors 789 
    -- successors 791 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_3993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_1_resize_ack_0, ack => cp_elements(790)); -- 
    scale_rename_req_3997_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(790), ack => array_obj_ref_1040_index_1_rename_req_0); -- 
    -- CP-element group 791 transition  input  no-bypass 
    -- predecessors 790 
    -- successors 784 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_3998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_1_rename_ack_0, ack => cp_elements(791)); -- 
    -- CP-element group 792 transition  input  output  no-bypass 
    -- predecessors 784 
    -- successors 793 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_sum_1_ack_0, ack => cp_elements(792)); -- 
    partial_sum_1_cr_4004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(792), ack => array_obj_ref_1040_index_sum_1_req_1); -- 
    -- CP-element group 793 transition  input  output  no-bypass 
    -- predecessors 792 
    -- successors 794 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_sum_1_ack_1, ack => cp_elements(793)); -- 
    final_index_req_4006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(793), ack => array_obj_ref_1040_offset_inst_req_0); -- 
    -- CP-element group 794 transition  input  output  no-bypass 
    -- predecessors 793 
    -- successors 795 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_offset_inst_ack_0, ack => cp_elements(794)); -- 
    sum_rename_req_4011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(794), ack => array_obj_ref_1040_root_address_inst_req_0); -- 
    -- CP-element group 795 transition  input  no-bypass 
    -- predecessors 794 
    -- successors 782 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1040_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_root_address_inst_ack_0, ack => cp_elements(795)); -- 
    -- CP-element group 796 transition  output  bypass 
    -- predecessors 782 
    -- successors 797 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1041_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1041_complete/final_reg_req
      -- 
    cp_elements(796) <= cp_elements(782);
    final_reg_req_4016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(796), ack => addr_of_1041_final_reg_req_0); -- 
    -- CP-element group 797 transition  input  no-bypass 
    -- predecessors 796 
    -- successors 783 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1041_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1041_complete/final_reg_ack
      -- 
    final_reg_ack_4017_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1041_final_reg_ack_0, ack => cp_elements(797)); -- 
    -- CP-element group 798 transition  bypass 
    -- predecessors 367 
    -- successors 799 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1047_trigger_
      -- 
    cp_elements(798) <= cp_elements(367);
    -- CP-element group 799 join  fork  transition  no-bypass 
    -- predecessors 798 812 
    -- successors 800 813 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1047_active_
      -- 
    cpelement_group_799 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(798);
      predecessors(1) <= cp_elements(812);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(799)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(799),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 800 join  transition  output  bypass 
    -- predecessors 799 814 
    -- successors 1125 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1047_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1048_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1048_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1048_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1180_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1180_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1180_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_addr_resize/base_resize_req
      -- 
    cpelement_group_800 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(799);
      predecessors(1) <= cp_elements(814);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(800)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(800),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5278_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(800), ack => ptr_deref_1181_base_resize_req_0); -- 
    -- CP-element group 801 join  transition  output  bypass 
    -- predecessors 805 808 
    -- successors 809 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_indices_scaled
      -- 
    cpelement_group_801 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(805);
      predecessors(1) <= cp_elements(808);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(801)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(801),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(801), ack => array_obj_ref_1046_index_sum_1_req_0); -- 
    -- CP-element group 802 transition  output  bypass 
    -- predecessors 724 
    -- successors 803 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1044_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1044_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1044_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_0/index_resize_req
      -- 
    cp_elements(802) <= cp_elements(724);
    index_resize_req_4035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(802), ack => array_obj_ref_1046_index_0_resize_req_0); -- 
    -- CP-element group 803 transition  input  output  no-bypass 
    -- predecessors 802 
    -- successors 804 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_0/scale_rr
      -- 
    index_resize_ack_4036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_0_resize_ack_0, ack => cp_elements(803)); -- 
    scale_rr_4040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(803), ack => array_obj_ref_1046_index_0_scale_req_0); -- 
    -- CP-element group 804 transition  input  output  no-bypass 
    -- predecessors 803 
    -- successors 805 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_0/scale_cr
      -- 
    scale_ra_4041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_0_scale_ack_0, ack => cp_elements(804)); -- 
    scale_cr_4042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(804), ack => array_obj_ref_1046_index_0_scale_req_1); -- 
    -- CP-element group 805 transition  input  no-bypass 
    -- predecessors 804 
    -- successors 801 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_0/scale_ca
      -- 
    scale_ca_4043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_0_scale_ack_1, ack => cp_elements(805)); -- 
    -- CP-element group 806 transition  output  bypass 
    -- predecessors 367 
    -- successors 807 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1045_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1045_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1045_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_1/$entry
      -- 
    cp_elements(806) <= cp_elements(367);
    index_resize_req_4052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(806), ack => array_obj_ref_1046_index_1_resize_req_0); -- 
    -- CP-element group 807 transition  input  output  no-bypass 
    -- predecessors 806 
    -- successors 808 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_resized_1
      -- 
    index_resize_ack_4053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_1_resize_ack_0, ack => cp_elements(807)); -- 
    scale_rename_req_4057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(807), ack => array_obj_ref_1046_index_1_rename_req_0); -- 
    -- CP-element group 808 transition  input  no-bypass 
    -- predecessors 807 
    -- successors 801 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_1_rename_ack_0, ack => cp_elements(808)); -- 
    -- CP-element group 809 transition  input  output  no-bypass 
    -- predecessors 801 
    -- successors 810 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_sum_1_ack_0, ack => cp_elements(809)); -- 
    partial_sum_1_cr_4064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(809), ack => array_obj_ref_1046_index_sum_1_req_1); -- 
    -- CP-element group 810 transition  input  output  no-bypass 
    -- predecessors 809 
    -- successors 811 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_sum_1_ack_1, ack => cp_elements(810)); -- 
    final_index_req_4066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(810), ack => array_obj_ref_1046_offset_inst_req_0); -- 
    -- CP-element group 811 transition  input  output  no-bypass 
    -- predecessors 810 
    -- successors 812 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_base_plus_offset/$entry
      -- 
    final_index_ack_4067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_offset_inst_ack_0, ack => cp_elements(811)); -- 
    sum_rename_req_4071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(811), ack => array_obj_ref_1046_root_address_inst_req_0); -- 
    -- CP-element group 812 transition  input  no-bypass 
    -- predecessors 811 
    -- successors 799 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1046_base_plus_offset/$exit
      -- 
    sum_rename_ack_4072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_root_address_inst_ack_0, ack => cp_elements(812)); -- 
    -- CP-element group 813 transition  output  bypass 
    -- predecessors 799 
    -- successors 814 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1047_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1047_complete/final_reg_req
      -- 
    cp_elements(813) <= cp_elements(799);
    final_reg_req_4076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(813), ack => addr_of_1047_final_reg_req_0); -- 
    -- CP-element group 814 transition  input  no-bypass 
    -- predecessors 813 
    -- successors 800 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1047_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1047_complete/final_reg_ack
      -- 
    final_reg_ack_4077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1047_final_reg_ack_0, ack => cp_elements(814)); -- 
    -- CP-element group 815 transition  bypass 
    -- predecessors 367 
    -- successors 816 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1053_trigger_
      -- 
    cp_elements(815) <= cp_elements(367);
    -- CP-element group 816 join  fork  transition  no-bypass 
    -- predecessors 815 829 
    -- successors 817 830 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1053_active_
      -- 
    cpelement_group_816 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(815);
      predecessors(1) <= cp_elements(829);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(816)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(816),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 817 join  transition  output  bypass 
    -- predecessors 816 831 
    -- successors 1115 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1054_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1054_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1054_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1053_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1176_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1176_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1176_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_addr_resize/base_resize_req
      -- 
    cpelement_group_817 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(816);
      predecessors(1) <= cp_elements(831);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(817)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(817),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(817), ack => ptr_deref_1177_base_resize_req_0); -- 
    -- CP-element group 818 join  transition  output  bypass 
    -- predecessors 822 825 
    -- successors 826 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/partial_sum_1_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/$entry
      -- 
    cpelement_group_818 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(822);
      predecessors(1) <= cp_elements(825);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(818)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(818),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4122_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(818), ack => array_obj_ref_1052_index_sum_1_req_0); -- 
    -- CP-element group 819 transition  output  bypass 
    -- predecessors 669 
    -- successors 820 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_0/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1050_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1050_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1050_active_
      -- 
    cp_elements(819) <= cp_elements(669);
    index_resize_req_4095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(819), ack => array_obj_ref_1052_index_0_resize_req_0); -- 
    -- CP-element group 820 transition  input  output  no-bypass 
    -- predecessors 819 
    -- successors 821 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_0/scale_rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_0/$exit
      -- 
    index_resize_ack_4096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_index_0_resize_ack_0, ack => cp_elements(820)); -- 
    scale_rr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(820), ack => array_obj_ref_1052_index_0_scale_req_0); -- 
    -- CP-element group 821 transition  input  output  no-bypass 
    -- predecessors 820 
    -- successors 822 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_0/scale_cr
      -- 
    scale_ra_4101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_index_0_scale_ack_0, ack => cp_elements(821)); -- 
    scale_cr_4102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(821), ack => array_obj_ref_1052_index_0_scale_req_1); -- 
    -- CP-element group 822 transition  input  no-bypass 
    -- predecessors 821 
    -- successors 818 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_0/scale_ca
      -- 
    scale_ca_4103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_index_0_scale_ack_1, ack => cp_elements(822)); -- 
    -- CP-element group 823 transition  output  bypass 
    -- predecessors 367 
    -- successors 824 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1051_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1051_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_1/index_resize_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1051_active_
      -- 
    cp_elements(823) <= cp_elements(367);
    index_resize_req_4112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(823), ack => array_obj_ref_1052_index_1_resize_req_0); -- 
    -- CP-element group 824 transition  input  output  no-bypass 
    -- predecessors 823 
    -- successors 825 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_1/scale_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_resize_1/$exit
      -- 
    index_resize_ack_4113_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_index_1_resize_ack_0, ack => cp_elements(824)); -- 
    scale_rename_req_4117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(824), ack => array_obj_ref_1052_index_1_rename_req_0); -- 
    -- CP-element group 825 transition  input  no-bypass 
    -- predecessors 824 
    -- successors 818 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_1/scale_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_index_scale_1/$exit
      -- 
    scale_rename_ack_4118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_index_1_rename_ack_0, ack => cp_elements(825)); -- 
    -- CP-element group 826 transition  input  output  no-bypass 
    -- predecessors 818 
    -- successors 827 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/partial_sum_1_cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/partial_sum_1_ra
      -- 
    partial_sum_1_ra_4123_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_index_sum_1_ack_0, ack => cp_elements(826)); -- 
    partial_sum_1_cr_4124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(826), ack => array_obj_ref_1052_index_sum_1_req_1); -- 
    -- CP-element group 827 transition  input  output  no-bypass 
    -- predecessors 826 
    -- successors 828 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4125_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_index_sum_1_ack_1, ack => cp_elements(827)); -- 
    final_index_req_4126_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(827), ack => array_obj_ref_1052_offset_inst_req_0); -- 
    -- CP-element group 828 transition  input  output  no-bypass 
    -- predecessors 827 
    -- successors 829 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4127_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_offset_inst_ack_0, ack => cp_elements(828)); -- 
    sum_rename_req_4131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => array_obj_ref_1052_root_address_inst_req_0); -- 
    -- CP-element group 829 transition  input  no-bypass 
    -- predecessors 828 
    -- successors 816 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1052_base_plus_offset/$exit
      -- 
    sum_rename_ack_4132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1052_root_address_inst_ack_0, ack => cp_elements(829)); -- 
    -- CP-element group 830 transition  output  bypass 
    -- predecessors 816 
    -- successors 831 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1053_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1053_complete/final_reg_req
      -- 
    cp_elements(830) <= cp_elements(816);
    final_reg_req_4136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(830), ack => addr_of_1053_final_reg_req_0); -- 
    -- CP-element group 831 transition  input  no-bypass 
    -- predecessors 830 
    -- successors 817 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1053_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1053_complete/final_reg_ack
      -- 
    final_reg_ack_4137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1053_final_reg_ack_0, ack => cp_elements(831)); -- 
    -- CP-element group 832 transition  bypass 
    -- predecessors 367 
    -- successors 833 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1059_trigger_
      -- 
    cp_elements(832) <= cp_elements(367);
    -- CP-element group 833 join  fork  transition  no-bypass 
    -- predecessors 832 846 
    -- successors 834 847 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1059_active_
      -- 
    cpelement_group_833 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(832);
      predecessors(1) <= cp_elements(846);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(833)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(833),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 834 join  transition  output  bypass 
    -- predecessors 833 848 
    -- successors 1250 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1060_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1060_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1060_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1059_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1244_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1244_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1244_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_addr_resize/base_resize_req
      -- 
    cpelement_group_834 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(833);
      predecessors(1) <= cp_elements(848);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(834)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(834),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(834), ack => ptr_deref_1245_base_resize_req_0); -- 
    -- CP-element group 835 join  transition  output  bypass 
    -- predecessors 839 842 
    -- successors 843 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_835 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(839);
      predecessors(1) <= cp_elements(842);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(835)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(835),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(835), ack => array_obj_ref_1058_index_sum_1_req_0); -- 
    -- CP-element group 836 transition  output  bypass 
    -- predecessors 676 
    -- successors 837 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1056_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1056_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1056_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_0/index_resize_req
      -- 
    cp_elements(836) <= cp_elements(676);
    index_resize_req_4155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(836), ack => array_obj_ref_1058_index_0_resize_req_0); -- 
    -- CP-element group 837 transition  input  output  no-bypass 
    -- predecessors 836 
    -- successors 838 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_0/scale_rr
      -- 
    index_resize_ack_4156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_0_resize_ack_0, ack => cp_elements(837)); -- 
    scale_rr_4160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(837), ack => array_obj_ref_1058_index_0_scale_req_0); -- 
    -- CP-element group 838 transition  input  output  no-bypass 
    -- predecessors 837 
    -- successors 839 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_0/scale_cr
      -- 
    scale_ra_4161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_0_scale_ack_0, ack => cp_elements(838)); -- 
    scale_cr_4162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(838), ack => array_obj_ref_1058_index_0_scale_req_1); -- 
    -- CP-element group 839 transition  input  no-bypass 
    -- predecessors 838 
    -- successors 835 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_0/scale_ca
      -- 
    scale_ca_4163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_0_scale_ack_1, ack => cp_elements(839)); -- 
    -- CP-element group 840 transition  output  bypass 
    -- predecessors 367 
    -- successors 841 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1057_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1057_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1057_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_1/index_resize_req
      -- 
    cp_elements(840) <= cp_elements(367);
    index_resize_req_4172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(840), ack => array_obj_ref_1058_index_1_resize_req_0); -- 
    -- CP-element group 841 transition  input  output  no-bypass 
    -- predecessors 840 
    -- successors 842 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_1_resize_ack_0, ack => cp_elements(841)); -- 
    scale_rename_req_4177_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(841), ack => array_obj_ref_1058_index_1_rename_req_0); -- 
    -- CP-element group 842 transition  input  no-bypass 
    -- predecessors 841 
    -- successors 835 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_1_rename_ack_0, ack => cp_elements(842)); -- 
    -- CP-element group 843 transition  input  output  no-bypass 
    -- predecessors 835 
    -- successors 844 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_sum_1_ack_0, ack => cp_elements(843)); -- 
    partial_sum_1_cr_4184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(843), ack => array_obj_ref_1058_index_sum_1_req_1); -- 
    -- CP-element group 844 transition  input  output  no-bypass 
    -- predecessors 843 
    -- successors 845 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_index_sum_1_ack_1, ack => cp_elements(844)); -- 
    final_index_req_4186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(844), ack => array_obj_ref_1058_offset_inst_req_0); -- 
    -- CP-element group 845 transition  input  output  no-bypass 
    -- predecessors 844 
    -- successors 846 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_offset_inst_ack_0, ack => cp_elements(845)); -- 
    sum_rename_req_4191_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(845), ack => array_obj_ref_1058_root_address_inst_req_0); -- 
    -- CP-element group 846 transition  input  no-bypass 
    -- predecessors 845 
    -- successors 833 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1058_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1058_root_address_inst_ack_0, ack => cp_elements(846)); -- 
    -- CP-element group 847 transition  output  bypass 
    -- predecessors 833 
    -- successors 848 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1059_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1059_complete/final_reg_req
      -- 
    cp_elements(847) <= cp_elements(833);
    final_reg_req_4196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(847), ack => addr_of_1059_final_reg_req_0); -- 
    -- CP-element group 848 transition  input  no-bypass 
    -- predecessors 847 
    -- successors 834 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1059_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1059_complete/final_reg_ack
      -- 
    final_reg_ack_4197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1059_final_reg_ack_0, ack => cp_elements(848)); -- 
    -- CP-element group 849 transition  bypass 
    -- predecessors 367 
    -- successors 850 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1065_trigger_
      -- 
    cp_elements(849) <= cp_elements(367);
    -- CP-element group 850 join  fork  transition  no-bypass 
    -- predecessors 849 863 
    -- successors 851 864 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1065_active_
      -- 
    cpelement_group_850 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(849);
      predecessors(1) <= cp_elements(863);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(850)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(850),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 851 join  transition  output  bypass 
    -- predecessors 850 865 
    -- successors 1240 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1066_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1066_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1066_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1065_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1240_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1240_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1240_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_addr_resize/base_resize_req
      -- 
    cpelement_group_851 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(850);
      predecessors(1) <= cp_elements(865);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(851)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(851),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(851), ack => ptr_deref_1241_base_resize_req_0); -- 
    -- CP-element group 852 join  transition  output  bypass 
    -- predecessors 856 859 
    -- successors 860 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_852 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(856);
      predecessors(1) <= cp_elements(859);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(852)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(852),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4242_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(852), ack => array_obj_ref_1064_index_sum_1_req_0); -- 
    -- CP-element group 853 transition  output  bypass 
    -- predecessors 700 
    -- successors 854 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1062_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1062_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1062_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_0/index_resize_req
      -- 
    cp_elements(853) <= cp_elements(700);
    index_resize_req_4215_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(853), ack => array_obj_ref_1064_index_0_resize_req_0); -- 
    -- CP-element group 854 transition  input  output  no-bypass 
    -- predecessors 853 
    -- successors 855 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_0/scale_rr
      -- 
    index_resize_ack_4216_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_index_0_resize_ack_0, ack => cp_elements(854)); -- 
    scale_rr_4220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(854), ack => array_obj_ref_1064_index_0_scale_req_0); -- 
    -- CP-element group 855 transition  input  output  no-bypass 
    -- predecessors 854 
    -- successors 856 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_0/scale_cr
      -- 
    scale_ra_4221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_index_0_scale_ack_0, ack => cp_elements(855)); -- 
    scale_cr_4222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(855), ack => array_obj_ref_1064_index_0_scale_req_1); -- 
    -- CP-element group 856 transition  input  no-bypass 
    -- predecessors 855 
    -- successors 852 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_0/scale_ca
      -- 
    scale_ca_4223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_index_0_scale_ack_1, ack => cp_elements(856)); -- 
    -- CP-element group 857 transition  output  bypass 
    -- predecessors 367 
    -- successors 858 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1063_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1063_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1063_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_1/index_resize_req
      -- 
    cp_elements(857) <= cp_elements(367);
    index_resize_req_4232_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(857), ack => array_obj_ref_1064_index_1_resize_req_0); -- 
    -- CP-element group 858 transition  input  output  no-bypass 
    -- predecessors 857 
    -- successors 859 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4233_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_index_1_resize_ack_0, ack => cp_elements(858)); -- 
    scale_rename_req_4237_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(858), ack => array_obj_ref_1064_index_1_rename_req_0); -- 
    -- CP-element group 859 transition  input  no-bypass 
    -- predecessors 858 
    -- successors 852 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_index_1_rename_ack_0, ack => cp_elements(859)); -- 
    -- CP-element group 860 transition  input  output  no-bypass 
    -- predecessors 852 
    -- successors 861 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4243_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_index_sum_1_ack_0, ack => cp_elements(860)); -- 
    partial_sum_1_cr_4244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(860), ack => array_obj_ref_1064_index_sum_1_req_1); -- 
    -- CP-element group 861 transition  input  output  no-bypass 
    -- predecessors 860 
    -- successors 862 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_index_sum_1_ack_1, ack => cp_elements(861)); -- 
    final_index_req_4246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(861), ack => array_obj_ref_1064_offset_inst_req_0); -- 
    -- CP-element group 862 transition  input  output  no-bypass 
    -- predecessors 861 
    -- successors 863 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_offset_inst_ack_0, ack => cp_elements(862)); -- 
    sum_rename_req_4251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(862), ack => array_obj_ref_1064_root_address_inst_req_0); -- 
    -- CP-element group 863 transition  input  no-bypass 
    -- predecessors 862 
    -- successors 850 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1064_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1064_root_address_inst_ack_0, ack => cp_elements(863)); -- 
    -- CP-element group 864 transition  output  bypass 
    -- predecessors 850 
    -- successors 865 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1065_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1065_complete/final_reg_req
      -- 
    cp_elements(864) <= cp_elements(850);
    final_reg_req_4256_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(864), ack => addr_of_1065_final_reg_req_0); -- 
    -- CP-element group 865 transition  input  no-bypass 
    -- predecessors 864 
    -- successors 851 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1065_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1065_complete/final_reg_ack
      -- 
    final_reg_ack_4257_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1065_final_reg_ack_0, ack => cp_elements(865)); -- 
    -- CP-element group 866 transition  bypass 
    -- predecessors 367 
    -- successors 867 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1071_trigger_
      -- 
    cp_elements(866) <= cp_elements(367);
    -- CP-element group 867 join  fork  transition  no-bypass 
    -- predecessors 866 880 
    -- successors 868 881 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1071_active_
      -- 
    cpelement_group_867 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(866);
      predecessors(1) <= cp_elements(880);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(867)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(867),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 868 join  transition  output  bypass 
    -- predecessors 867 882 
    -- successors 1230 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1072_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1072_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1072_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1071_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1236_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1236_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1236_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_addr_resize/base_resize_req
      -- 
    cpelement_group_868 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(867);
      predecessors(1) <= cp_elements(882);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(868)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(868),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5662_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => ptr_deref_1237_base_resize_req_0); -- 
    -- CP-element group 869 join  transition  output  bypass 
    -- predecessors 873 876 
    -- successors 877 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_869 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(873);
      predecessors(1) <= cp_elements(876);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(869)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(869),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(869), ack => array_obj_ref_1070_index_sum_1_req_0); -- 
    -- CP-element group 870 transition  output  bypass 
    -- predecessors 724 
    -- successors 871 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1068_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1068_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1068_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_0/index_resize_req
      -- 
    cp_elements(870) <= cp_elements(724);
    index_resize_req_4275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(870), ack => array_obj_ref_1070_index_0_resize_req_0); -- 
    -- CP-element group 871 transition  input  output  no-bypass 
    -- predecessors 870 
    -- successors 872 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_0/scale_rr
      -- 
    index_resize_ack_4276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_index_0_resize_ack_0, ack => cp_elements(871)); -- 
    scale_rr_4280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(871), ack => array_obj_ref_1070_index_0_scale_req_0); -- 
    -- CP-element group 872 transition  input  output  no-bypass 
    -- predecessors 871 
    -- successors 873 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_0/scale_cr
      -- 
    scale_ra_4281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_index_0_scale_ack_0, ack => cp_elements(872)); -- 
    scale_cr_4282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(872), ack => array_obj_ref_1070_index_0_scale_req_1); -- 
    -- CP-element group 873 transition  input  no-bypass 
    -- predecessors 872 
    -- successors 869 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_0/scale_ca
      -- 
    scale_ca_4283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_index_0_scale_ack_1, ack => cp_elements(873)); -- 
    -- CP-element group 874 transition  output  bypass 
    -- predecessors 367 
    -- successors 875 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1069_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1069_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1069_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_1/index_resize_req
      -- 
    cp_elements(874) <= cp_elements(367);
    index_resize_req_4292_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(874), ack => array_obj_ref_1070_index_1_resize_req_0); -- 
    -- CP-element group 875 transition  input  output  no-bypass 
    -- predecessors 874 
    -- successors 876 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4293_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_index_1_resize_ack_0, ack => cp_elements(875)); -- 
    scale_rename_req_4297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(875), ack => array_obj_ref_1070_index_1_rename_req_0); -- 
    -- CP-element group 876 transition  input  no-bypass 
    -- predecessors 875 
    -- successors 869 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_index_1_rename_ack_0, ack => cp_elements(876)); -- 
    -- CP-element group 877 transition  input  output  no-bypass 
    -- predecessors 869 
    -- successors 878 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_index_sum_1_ack_0, ack => cp_elements(877)); -- 
    partial_sum_1_cr_4304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(877), ack => array_obj_ref_1070_index_sum_1_req_1); -- 
    -- CP-element group 878 transition  input  output  no-bypass 
    -- predecessors 877 
    -- successors 879 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_index_sum_1_ack_1, ack => cp_elements(878)); -- 
    final_index_req_4306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(878), ack => array_obj_ref_1070_offset_inst_req_0); -- 
    -- CP-element group 879 transition  input  output  no-bypass 
    -- predecessors 878 
    -- successors 880 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_offset_inst_ack_0, ack => cp_elements(879)); -- 
    sum_rename_req_4311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(879), ack => array_obj_ref_1070_root_address_inst_req_0); -- 
    -- CP-element group 880 transition  input  no-bypass 
    -- predecessors 879 
    -- successors 867 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1070_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1070_root_address_inst_ack_0, ack => cp_elements(880)); -- 
    -- CP-element group 881 transition  output  bypass 
    -- predecessors 867 
    -- successors 882 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1071_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1071_complete/final_reg_req
      -- 
    cp_elements(881) <= cp_elements(867);
    final_reg_req_4316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(881), ack => addr_of_1071_final_reg_req_0); -- 
    -- CP-element group 882 transition  input  no-bypass 
    -- predecessors 881 
    -- successors 868 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1071_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1071_complete/final_reg_ack
      -- 
    final_reg_ack_4317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1071_final_reg_ack_0, ack => cp_elements(882)); -- 
    -- CP-element group 883 transition  bypass 
    -- predecessors 367 
    -- successors 884 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1077_trigger_
      -- 
    cp_elements(883) <= cp_elements(367);
    -- CP-element group 884 join  fork  transition  no-bypass 
    -- predecessors 883 897 
    -- successors 885 898 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1077_active_
      -- 
    cpelement_group_884 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(883);
      predecessors(1) <= cp_elements(897);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(884)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(884),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 885 join  transition  output  bypass 
    -- predecessors 884 899 
    -- successors 1220 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1078_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1078_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1078_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1077_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1232_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1232_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1232_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_addr_resize/base_resize_req
      -- 
    cpelement_group_885 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(884);
      predecessors(1) <= cp_elements(899);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(885)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(885),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(885), ack => ptr_deref_1233_base_resize_req_0); -- 
    -- CP-element group 886 join  transition  output  bypass 
    -- predecessors 890 893 
    -- successors 894 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_886 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(890);
      predecessors(1) <= cp_elements(893);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(886)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(886),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4362_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(886), ack => array_obj_ref_1076_index_sum_1_req_0); -- 
    -- CP-element group 887 transition  output  bypass 
    -- predecessors 669 
    -- successors 888 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1074_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1074_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1074_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_0/index_resize_req
      -- 
    cp_elements(887) <= cp_elements(669);
    index_resize_req_4335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(887), ack => array_obj_ref_1076_index_0_resize_req_0); -- 
    -- CP-element group 888 transition  input  output  no-bypass 
    -- predecessors 887 
    -- successors 889 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_0/scale_rr
      -- 
    index_resize_ack_4336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_index_0_resize_ack_0, ack => cp_elements(888)); -- 
    scale_rr_4340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(888), ack => array_obj_ref_1076_index_0_scale_req_0); -- 
    -- CP-element group 889 transition  input  output  no-bypass 
    -- predecessors 888 
    -- successors 890 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_0/scale_cr
      -- 
    scale_ra_4341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_index_0_scale_ack_0, ack => cp_elements(889)); -- 
    scale_cr_4342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(889), ack => array_obj_ref_1076_index_0_scale_req_1); -- 
    -- CP-element group 890 transition  input  no-bypass 
    -- predecessors 889 
    -- successors 886 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_0/scale_ca
      -- 
    scale_ca_4343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_index_0_scale_ack_1, ack => cp_elements(890)); -- 
    -- CP-element group 891 transition  output  bypass 
    -- predecessors 367 
    -- successors 892 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1075_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1075_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1075_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_1/index_resize_req
      -- 
    cp_elements(891) <= cp_elements(367);
    index_resize_req_4352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(891), ack => array_obj_ref_1076_index_1_resize_req_0); -- 
    -- CP-element group 892 transition  input  output  no-bypass 
    -- predecessors 891 
    -- successors 893 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_index_1_resize_ack_0, ack => cp_elements(892)); -- 
    scale_rename_req_4357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(892), ack => array_obj_ref_1076_index_1_rename_req_0); -- 
    -- CP-element group 893 transition  input  no-bypass 
    -- predecessors 892 
    -- successors 886 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_index_1_rename_ack_0, ack => cp_elements(893)); -- 
    -- CP-element group 894 transition  input  output  no-bypass 
    -- predecessors 886 
    -- successors 895 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_index_sum_1_ack_0, ack => cp_elements(894)); -- 
    partial_sum_1_cr_4364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(894), ack => array_obj_ref_1076_index_sum_1_req_1); -- 
    -- CP-element group 895 transition  input  output  no-bypass 
    -- predecessors 894 
    -- successors 896 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_index_sum_1_ack_1, ack => cp_elements(895)); -- 
    final_index_req_4366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(895), ack => array_obj_ref_1076_offset_inst_req_0); -- 
    -- CP-element group 896 transition  input  output  no-bypass 
    -- predecessors 895 
    -- successors 897 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4367_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_offset_inst_ack_0, ack => cp_elements(896)); -- 
    sum_rename_req_4371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(896), ack => array_obj_ref_1076_root_address_inst_req_0); -- 
    -- CP-element group 897 transition  input  no-bypass 
    -- predecessors 896 
    -- successors 884 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1076_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1076_root_address_inst_ack_0, ack => cp_elements(897)); -- 
    -- CP-element group 898 transition  output  bypass 
    -- predecessors 884 
    -- successors 899 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1077_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1077_complete/final_reg_req
      -- 
    cp_elements(898) <= cp_elements(884);
    final_reg_req_4376_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(898), ack => addr_of_1077_final_reg_req_0); -- 
    -- CP-element group 899 transition  input  no-bypass 
    -- predecessors 898 
    -- successors 885 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1077_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1077_complete/final_reg_ack
      -- 
    final_reg_ack_4377_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1077_final_reg_ack_0, ack => cp_elements(899)); -- 
    -- CP-element group 900 transition  bypass 
    -- predecessors 367 
    -- successors 901 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1083_trigger_
      -- 
    cp_elements(900) <= cp_elements(367);
    -- CP-element group 901 join  fork  transition  no-bypass 
    -- predecessors 900 914 
    -- successors 902 915 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1083_active_
      -- 
    cpelement_group_901 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(900);
      predecessors(1) <= cp_elements(914);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(901)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(901),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 902 join  transition  output  bypass 
    -- predecessors 901 916 
    -- successors 1355 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1084_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1084_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1084_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1083_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1300_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1300_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1300_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_addr_resize/base_resize_req
      -- 
    cpelement_group_902 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(901);
      predecessors(1) <= cp_elements(916);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(902)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(902),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_6150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(902), ack => ptr_deref_1301_base_resize_req_0); -- 
    -- CP-element group 903 join  transition  output  bypass 
    -- predecessors 907 910 
    -- successors 911 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_903 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(907);
      predecessors(1) <= cp_elements(910);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(903)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(903),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4422_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(903), ack => array_obj_ref_1082_index_sum_1_req_0); -- 
    -- CP-element group 904 transition  output  bypass 
    -- predecessors 676 
    -- successors 905 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1080_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1080_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1080_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_0/index_resize_req
      -- 
    cp_elements(904) <= cp_elements(676);
    index_resize_req_4395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(904), ack => array_obj_ref_1082_index_0_resize_req_0); -- 
    -- CP-element group 905 transition  input  output  no-bypass 
    -- predecessors 904 
    -- successors 906 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_0/scale_rr
      -- 
    index_resize_ack_4396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_index_0_resize_ack_0, ack => cp_elements(905)); -- 
    scale_rr_4400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(905), ack => array_obj_ref_1082_index_0_scale_req_0); -- 
    -- CP-element group 906 transition  input  output  no-bypass 
    -- predecessors 905 
    -- successors 907 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_0/scale_cr
      -- 
    scale_ra_4401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_index_0_scale_ack_0, ack => cp_elements(906)); -- 
    scale_cr_4402_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(906), ack => array_obj_ref_1082_index_0_scale_req_1); -- 
    -- CP-element group 907 transition  input  no-bypass 
    -- predecessors 906 
    -- successors 903 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_0/scale_ca
      -- 
    scale_ca_4403_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_index_0_scale_ack_1, ack => cp_elements(907)); -- 
    -- CP-element group 908 transition  output  bypass 
    -- predecessors 367 
    -- successors 909 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1081_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1081_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1081_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_1/index_resize_req
      -- 
    cp_elements(908) <= cp_elements(367);
    index_resize_req_4412_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(908), ack => array_obj_ref_1082_index_1_resize_req_0); -- 
    -- CP-element group 909 transition  input  output  no-bypass 
    -- predecessors 908 
    -- successors 910 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_index_1_resize_ack_0, ack => cp_elements(909)); -- 
    scale_rename_req_4417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(909), ack => array_obj_ref_1082_index_1_rename_req_0); -- 
    -- CP-element group 910 transition  input  no-bypass 
    -- predecessors 909 
    -- successors 903 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_index_1_rename_ack_0, ack => cp_elements(910)); -- 
    -- CP-element group 911 transition  input  output  no-bypass 
    -- predecessors 903 
    -- successors 912 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4423_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_index_sum_1_ack_0, ack => cp_elements(911)); -- 
    partial_sum_1_cr_4424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(911), ack => array_obj_ref_1082_index_sum_1_req_1); -- 
    -- CP-element group 912 transition  input  output  no-bypass 
    -- predecessors 911 
    -- successors 913 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_index_sum_1_ack_1, ack => cp_elements(912)); -- 
    final_index_req_4426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(912), ack => array_obj_ref_1082_offset_inst_req_0); -- 
    -- CP-element group 913 transition  input  output  no-bypass 
    -- predecessors 912 
    -- successors 914 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_offset_inst_ack_0, ack => cp_elements(913)); -- 
    sum_rename_req_4431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(913), ack => array_obj_ref_1082_root_address_inst_req_0); -- 
    -- CP-element group 914 transition  input  no-bypass 
    -- predecessors 913 
    -- successors 901 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1082_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1082_root_address_inst_ack_0, ack => cp_elements(914)); -- 
    -- CP-element group 915 transition  output  bypass 
    -- predecessors 901 
    -- successors 916 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1083_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1083_complete/final_reg_req
      -- 
    cp_elements(915) <= cp_elements(901);
    final_reg_req_4436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(915), ack => addr_of_1083_final_reg_req_0); -- 
    -- CP-element group 916 transition  input  no-bypass 
    -- predecessors 915 
    -- successors 902 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1083_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1083_complete/final_reg_ack
      -- 
    final_reg_ack_4437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1083_final_reg_ack_0, ack => cp_elements(916)); -- 
    -- CP-element group 917 transition  bypass 
    -- predecessors 367 
    -- successors 918 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1089_trigger_
      -- 
    cp_elements(917) <= cp_elements(367);
    -- CP-element group 918 join  fork  transition  no-bypass 
    -- predecessors 917 931 
    -- successors 919 932 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1089_active_
      -- 
    cpelement_group_918 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(917);
      predecessors(1) <= cp_elements(931);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(918)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(918),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 919 join  transition  output  bypass 
    -- predecessors 918 933 
    -- successors 1345 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1090_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1090_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1090_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1089_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1296_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1296_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1296_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_addr_resize/base_resize_req
      -- 
    cpelement_group_919 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(918);
      predecessors(1) <= cp_elements(933);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(919)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(919),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_6098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(919), ack => ptr_deref_1297_base_resize_req_0); -- 
    -- CP-element group 920 join  transition  output  bypass 
    -- predecessors 924 927 
    -- successors 928 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_920 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(924);
      predecessors(1) <= cp_elements(927);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(920)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(920),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(920), ack => array_obj_ref_1088_index_sum_1_req_0); -- 
    -- CP-element group 921 transition  output  bypass 
    -- predecessors 700 
    -- successors 922 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1086_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1086_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1086_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_0/index_resize_req
      -- 
    cp_elements(921) <= cp_elements(700);
    index_resize_req_4455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(921), ack => array_obj_ref_1088_index_0_resize_req_0); -- 
    -- CP-element group 922 transition  input  output  no-bypass 
    -- predecessors 921 
    -- successors 923 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_0/scale_rr
      -- 
    index_resize_ack_4456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_0_resize_ack_0, ack => cp_elements(922)); -- 
    scale_rr_4460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(922), ack => array_obj_ref_1088_index_0_scale_req_0); -- 
    -- CP-element group 923 transition  input  output  no-bypass 
    -- predecessors 922 
    -- successors 924 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_0/scale_cr
      -- 
    scale_ra_4461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_0_scale_ack_0, ack => cp_elements(923)); -- 
    scale_cr_4462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(923), ack => array_obj_ref_1088_index_0_scale_req_1); -- 
    -- CP-element group 924 transition  input  no-bypass 
    -- predecessors 923 
    -- successors 920 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_0/scale_ca
      -- 
    scale_ca_4463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_0_scale_ack_1, ack => cp_elements(924)); -- 
    -- CP-element group 925 transition  output  bypass 
    -- predecessors 367 
    -- successors 926 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1087_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1087_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1087_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_1/index_resize_req
      -- 
    cp_elements(925) <= cp_elements(367);
    index_resize_req_4472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(925), ack => array_obj_ref_1088_index_1_resize_req_0); -- 
    -- CP-element group 926 transition  input  output  no-bypass 
    -- predecessors 925 
    -- successors 927 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_1_resize_ack_0, ack => cp_elements(926)); -- 
    scale_rename_req_4477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(926), ack => array_obj_ref_1088_index_1_rename_req_0); -- 
    -- CP-element group 927 transition  input  no-bypass 
    -- predecessors 926 
    -- successors 920 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_1_rename_ack_0, ack => cp_elements(927)); -- 
    -- CP-element group 928 transition  input  output  no-bypass 
    -- predecessors 920 
    -- successors 929 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_sum_1_ack_0, ack => cp_elements(928)); -- 
    partial_sum_1_cr_4484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(928), ack => array_obj_ref_1088_index_sum_1_req_1); -- 
    -- CP-element group 929 transition  input  output  no-bypass 
    -- predecessors 928 
    -- successors 930 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_index_sum_1_ack_1, ack => cp_elements(929)); -- 
    final_index_req_4486_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(929), ack => array_obj_ref_1088_offset_inst_req_0); -- 
    -- CP-element group 930 transition  input  output  no-bypass 
    -- predecessors 929 
    -- successors 931 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4487_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_offset_inst_ack_0, ack => cp_elements(930)); -- 
    sum_rename_req_4491_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(930), ack => array_obj_ref_1088_root_address_inst_req_0); -- 
    -- CP-element group 931 transition  input  no-bypass 
    -- predecessors 930 
    -- successors 918 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1088_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4492_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1088_root_address_inst_ack_0, ack => cp_elements(931)); -- 
    -- CP-element group 932 transition  output  bypass 
    -- predecessors 918 
    -- successors 933 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1089_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1089_complete/final_reg_req
      -- 
    cp_elements(932) <= cp_elements(918);
    final_reg_req_4496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(932), ack => addr_of_1089_final_reg_req_0); -- 
    -- CP-element group 933 transition  input  no-bypass 
    -- predecessors 932 
    -- successors 919 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1089_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1089_complete/final_reg_ack
      -- 
    final_reg_ack_4497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1089_final_reg_ack_0, ack => cp_elements(933)); -- 
    -- CP-element group 934 transition  bypass 
    -- predecessors 367 
    -- successors 935 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1095_trigger_
      -- 
    cp_elements(934) <= cp_elements(367);
    -- CP-element group 935 join  fork  transition  no-bypass 
    -- predecessors 934 948 
    -- successors 936 949 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1095_active_
      -- 
    cpelement_group_935 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(934);
      predecessors(1) <= cp_elements(948);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(935)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(935),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 936 join  transition  output  bypass 
    -- predecessors 935 950 
    -- successors 1335 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1096_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1096_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1096_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1095_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1292_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1292_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1292_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_addr_resize/base_resize_req
      -- 
    cpelement_group_936 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(935);
      predecessors(1) <= cp_elements(950);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(936)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(936),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_6046_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(936), ack => ptr_deref_1293_base_resize_req_0); -- 
    -- CP-element group 937 join  transition  output  bypass 
    -- predecessors 941 944 
    -- successors 945 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_937 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(941);
      predecessors(1) <= cp_elements(944);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(937)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(937),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4542_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(937), ack => array_obj_ref_1094_index_sum_1_req_0); -- 
    -- CP-element group 938 transition  output  bypass 
    -- predecessors 724 
    -- successors 939 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1092_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1092_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1092_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_0/index_resize_req
      -- 
    cp_elements(938) <= cp_elements(724);
    index_resize_req_4515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(938), ack => array_obj_ref_1094_index_0_resize_req_0); -- 
    -- CP-element group 939 transition  input  output  no-bypass 
    -- predecessors 938 
    -- successors 940 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_0/scale_rr
      -- 
    index_resize_ack_4516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_index_0_resize_ack_0, ack => cp_elements(939)); -- 
    scale_rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => array_obj_ref_1094_index_0_scale_req_0); -- 
    -- CP-element group 940 transition  input  output  no-bypass 
    -- predecessors 939 
    -- successors 941 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_0/scale_cr
      -- 
    scale_ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_index_0_scale_ack_0, ack => cp_elements(940)); -- 
    scale_cr_4522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(940), ack => array_obj_ref_1094_index_0_scale_req_1); -- 
    -- CP-element group 941 transition  input  no-bypass 
    -- predecessors 940 
    -- successors 937 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_0/scale_ca
      -- 
    scale_ca_4523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_index_0_scale_ack_1, ack => cp_elements(941)); -- 
    -- CP-element group 942 transition  output  bypass 
    -- predecessors 367 
    -- successors 943 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1093_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1093_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1093_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_1/index_resize_req
      -- 
    cp_elements(942) <= cp_elements(367);
    index_resize_req_4532_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(942), ack => array_obj_ref_1094_index_1_resize_req_0); -- 
    -- CP-element group 943 transition  input  output  no-bypass 
    -- predecessors 942 
    -- successors 944 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_index_1_resize_ack_0, ack => cp_elements(943)); -- 
    scale_rename_req_4537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(943), ack => array_obj_ref_1094_index_1_rename_req_0); -- 
    -- CP-element group 944 transition  input  no-bypass 
    -- predecessors 943 
    -- successors 937 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4538_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_index_1_rename_ack_0, ack => cp_elements(944)); -- 
    -- CP-element group 945 transition  input  output  no-bypass 
    -- predecessors 937 
    -- successors 946 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4543_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_index_sum_1_ack_0, ack => cp_elements(945)); -- 
    partial_sum_1_cr_4544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(945), ack => array_obj_ref_1094_index_sum_1_req_1); -- 
    -- CP-element group 946 transition  input  output  no-bypass 
    -- predecessors 945 
    -- successors 947 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_index_sum_1_ack_1, ack => cp_elements(946)); -- 
    final_index_req_4546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(946), ack => array_obj_ref_1094_offset_inst_req_0); -- 
    -- CP-element group 947 transition  input  output  no-bypass 
    -- predecessors 946 
    -- successors 948 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_offset_inst_ack_0, ack => cp_elements(947)); -- 
    sum_rename_req_4551_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(947), ack => array_obj_ref_1094_root_address_inst_req_0); -- 
    -- CP-element group 948 transition  input  no-bypass 
    -- predecessors 947 
    -- successors 935 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1094_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4552_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1094_root_address_inst_ack_0, ack => cp_elements(948)); -- 
    -- CP-element group 949 transition  output  bypass 
    -- predecessors 935 
    -- successors 950 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1095_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1095_complete/final_reg_req
      -- 
    cp_elements(949) <= cp_elements(935);
    final_reg_req_4556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(949), ack => addr_of_1095_final_reg_req_0); -- 
    -- CP-element group 950 transition  input  no-bypass 
    -- predecessors 949 
    -- successors 936 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1095_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1095_complete/final_reg_ack
      -- 
    final_reg_ack_4557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1095_final_reg_ack_0, ack => cp_elements(950)); -- 
    -- CP-element group 951 transition  bypass 
    -- predecessors 367 
    -- successors 952 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1101_trigger_
      -- 
    cp_elements(951) <= cp_elements(367);
    -- CP-element group 952 join  fork  transition  no-bypass 
    -- predecessors 951 965 
    -- successors 953 966 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1101_active_
      -- 
    cpelement_group_952 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(951);
      predecessors(1) <= cp_elements(965);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(952)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(952),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 953 join  transition  output  bypass 
    -- predecessors 952 967 
    -- successors 1325 
    -- members (10) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1288_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1288_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1288_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1102_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1102_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1102_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1101_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_addr_resize/base_resize_req
      -- 
    cpelement_group_953 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(952);
      predecessors(1) <= cp_elements(967);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(953)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(953),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    base_resize_req_5994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(953), ack => ptr_deref_1289_base_resize_req_0); -- 
    -- CP-element group 954 join  transition  output  bypass 
    -- predecessors 958 961 
    -- successors 962 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_indices_scaled
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/partial_sum_1_rr
      -- 
    cpelement_group_954 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(958);
      predecessors(1) <= cp_elements(961);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(954)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(954),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    partial_sum_1_rr_4602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(954), ack => array_obj_ref_1100_index_sum_1_req_0); -- 
    -- CP-element group 955 transition  output  bypass 
    -- predecessors 669 
    -- successors 956 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_computed_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1098_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1098_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1098_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_0/index_resize_req
      -- 
    cp_elements(955) <= cp_elements(669);
    index_resize_req_4575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(955), ack => array_obj_ref_1100_index_0_resize_req_0); -- 
    -- CP-element group 956 transition  input  output  no-bypass 
    -- predecessors 955 
    -- successors 957 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resized_0
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_0/scale_rr
      -- 
    index_resize_ack_4576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_index_0_resize_ack_0, ack => cp_elements(956)); -- 
    scale_rr_4580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(956), ack => array_obj_ref_1100_index_0_scale_req_0); -- 
    -- CP-element group 957 transition  input  output  no-bypass 
    -- predecessors 956 
    -- successors 958 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_0/scale_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_0/scale_cr
      -- 
    scale_ra_4581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_index_0_scale_ack_0, ack => cp_elements(957)); -- 
    scale_cr_4582_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(957), ack => array_obj_ref_1100_index_0_scale_req_1); -- 
    -- CP-element group 958 transition  input  no-bypass 
    -- predecessors 957 
    -- successors 954 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_0/scale_ca
      -- 
    scale_ca_4583_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_index_0_scale_ack_1, ack => cp_elements(958)); -- 
    -- CP-element group 959 transition  output  bypass 
    -- predecessors 367 
    -- successors 960 
    -- members (6) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_computed_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1099_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1099_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1099_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_1/index_resize_req
      -- 
    cp_elements(959) <= cp_elements(367);
    index_resize_req_4592_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(959), ack => array_obj_ref_1100_index_1_resize_req_0); -- 
    -- CP-element group 960 transition  input  output  no-bypass 
    -- predecessors 959 
    -- successors 961 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resized_1
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_resize_1/index_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_1/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_1/scale_rename_req
      -- 
    index_resize_ack_4593_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_index_1_resize_ack_0, ack => cp_elements(960)); -- 
    scale_rename_req_4597_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(960), ack => array_obj_ref_1100_index_1_rename_req_0); -- 
    -- CP-element group 961 transition  input  no-bypass 
    -- predecessors 960 
    -- successors 954 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_1/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_index_scale_1/scale_rename_ack
      -- 
    scale_rename_ack_4598_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_index_1_rename_ack_0, ack => cp_elements(961)); -- 
    -- CP-element group 962 transition  input  output  no-bypass 
    -- predecessors 954 
    -- successors 963 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/partial_sum_1_ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/partial_sum_1_cr
      -- 
    partial_sum_1_ra_4603_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_index_sum_1_ack_0, ack => cp_elements(962)); -- 
    partial_sum_1_cr_4604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(962), ack => array_obj_ref_1100_index_sum_1_req_1); -- 
    -- CP-element group 963 transition  input  output  no-bypass 
    -- predecessors 962 
    -- successors 964 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/partial_sum_1_ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/final_index_req
      -- 
    partial_sum_1_ca_4605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_index_sum_1_ack_1, ack => cp_elements(963)); -- 
    final_index_req_4606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(963), ack => array_obj_ref_1100_offset_inst_req_0); -- 
    -- CP-element group 964 transition  input  output  no-bypass 
    -- predecessors 963 
    -- successors 965 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_offset_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_add_indices/final_index_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_offset_inst_ack_0, ack => cp_elements(964)); -- 
    sum_rename_req_4611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(964), ack => array_obj_ref_1100_root_address_inst_req_0); -- 
    -- CP-element group 965 transition  input  no-bypass 
    -- predecessors 964 
    -- successors 952 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/array_obj_ref_1100_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1100_root_address_inst_ack_0, ack => cp_elements(965)); -- 
    -- CP-element group 966 transition  output  bypass 
    -- predecessors 952 
    -- successors 967 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1101_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1101_complete/final_reg_req
      -- 
    cp_elements(966) <= cp_elements(952);
    final_reg_req_4616_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(966), ack => addr_of_1101_final_reg_req_0); -- 
    -- CP-element group 967 transition  input  no-bypass 
    -- predecessors 966 
    -- successors 953 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1101_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/addr_of_1101_complete/final_reg_ack
      -- 
    final_reg_ack_4617_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1101_final_reg_ack_0, ack => cp_elements(967)); -- 
    -- CP-element group 968 join  fork  transition  bypass 
    -- predecessors 972 974 
    -- successors 969 975 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_active_
      -- 
    cpelement_group_968 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(972);
      predecessors(1) <= cp_elements(974);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(968)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(968),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 969 join  fork  transition  bypass 
    -- predecessors 968 977 
    -- successors 1051 1156 1261 1366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1106_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1106_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1106_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_completed_
      -- 
    cpelement_group_969 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(968);
      predecessors(1) <= cp_elements(977);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(969)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(969),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 970 transition  input  output  no-bypass 
    -- predecessors 377 
    -- successors 971 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_base_resize_ack_0, ack => cp_elements(970)); -- 
    sum_rename_req_4639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(970), ack => ptr_deref_1105_root_address_inst_req_0); -- 
    -- CP-element group 971 transition  input  output  no-bypass 
    -- predecessors 970 
    -- successors 972 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_root_address_inst_ack_0, ack => cp_elements(971)); -- 
    root_register_req_4644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(971), ack => ptr_deref_1105_addr_0_req_0); -- 
    -- CP-element group 972 fork  transition  input  no-bypass 
    -- predecessors 971 
    -- successors 968 973 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_word_addrgen/root_register_ack
      -- 
    root_register_ack_4645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_addr_0_ack_0, ack => cp_elements(972)); -- 
    -- CP-element group 973 transition  output  bypass 
    -- predecessors 972 
    -- successors 974 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/word_access/word_access_0/rr
      -- 
    cp_elements(973) <= cp_elements(972);
    rr_4655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(973), ack => ptr_deref_1105_load_0_req_0); -- 
    -- CP-element group 974 transition  input  no-bypass 
    -- predecessors 973 
    -- successors 968 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_request/word_access/word_access_0/ra
      -- 
    ra_4656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_load_0_ack_0, ack => cp_elements(974)); -- 
    -- CP-element group 975 transition  output  bypass 
    -- predecessors 968 
    -- successors 976 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/word_access/word_access_0/cr
      -- 
    cp_elements(975) <= cp_elements(968);
    cr_4666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(975), ack => ptr_deref_1105_load_0_req_1); -- 
    -- CP-element group 976 transition  input  output  no-bypass 
    -- predecessors 975 
    -- successors 977 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/merge_req
      -- 
    ca_4667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_load_0_ack_1, ack => cp_elements(976)); -- 
    merge_req_4668_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(976), ack => ptr_deref_1105_gather_scatter_req_0); -- 
    -- CP-element group 977 transition  input  no-bypass 
    -- predecessors 976 
    -- successors 969 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1105_complete/merge_ack
      -- 
    merge_ack_4669_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_gather_scatter_ack_0, ack => cp_elements(977)); -- 
    -- CP-element group 978 join  fork  transition  bypass 
    -- predecessors 982 984 
    -- successors 979 985 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_active_
      -- 
    cpelement_group_978 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(982);
      predecessors(1) <= cp_elements(984);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(978)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(978),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 979 join  fork  transition  bypass 
    -- predecessors 978 987 
    -- successors 1052 1472 1772 2072 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1110_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1110_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1110_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_completed_
      -- 
    cpelement_group_979 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(978);
      predecessors(1) <= cp_elements(987);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(979)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(979),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 980 transition  input  output  no-bypass 
    -- predecessors 749 
    -- successors 981 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4687_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_base_resize_ack_0, ack => cp_elements(980)); -- 
    sum_rename_req_4691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(980), ack => ptr_deref_1109_root_address_inst_req_0); -- 
    -- CP-element group 981 transition  input  output  no-bypass 
    -- predecessors 980 
    -- successors 982 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_root_address_inst_ack_0, ack => cp_elements(981)); -- 
    root_register_req_4696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(981), ack => ptr_deref_1109_addr_0_req_0); -- 
    -- CP-element group 982 fork  transition  input  no-bypass 
    -- predecessors 981 
    -- successors 978 983 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_word_addrgen/root_register_ack
      -- 
    root_register_ack_4697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_addr_0_ack_0, ack => cp_elements(982)); -- 
    -- CP-element group 983 transition  output  bypass 
    -- predecessors 982 
    -- successors 984 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/word_access/word_access_0/rr
      -- 
    cp_elements(983) <= cp_elements(982);
    rr_4707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(983), ack => ptr_deref_1109_load_0_req_0); -- 
    -- CP-element group 984 transition  input  no-bypass 
    -- predecessors 983 
    -- successors 978 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_request/word_access/word_access_0/ra
      -- 
    ra_4708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_load_0_ack_0, ack => cp_elements(984)); -- 
    -- CP-element group 985 transition  output  bypass 
    -- predecessors 978 
    -- successors 986 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/word_access/word_access_0/cr
      -- 
    cp_elements(985) <= cp_elements(978);
    cr_4718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(985), ack => ptr_deref_1109_load_0_req_1); -- 
    -- CP-element group 986 transition  input  output  no-bypass 
    -- predecessors 985 
    -- successors 987 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/merge_req
      -- 
    ca_4719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_load_0_ack_1, ack => cp_elements(986)); -- 
    merge_req_4720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(986), ack => ptr_deref_1109_gather_scatter_req_0); -- 
    -- CP-element group 987 transition  input  no-bypass 
    -- predecessors 986 
    -- successors 979 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1109_complete/merge_ack
      -- 
    merge_ack_4721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_gather_scatter_ack_0, ack => cp_elements(987)); -- 
    -- CP-element group 988 join  fork  transition  bypass 
    -- predecessors 992 994 
    -- successors 989 995 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_active_
      -- 
    cpelement_group_988 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(992);
      predecessors(1) <= cp_elements(994);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(988)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(988),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 989 join  fork  transition  bypass 
    -- predecessors 988 997 
    -- successors 1060 1165 1270 1375 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1114_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1114_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1114_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_completed_
      -- 
    cpelement_group_989 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(988);
      predecessors(1) <= cp_elements(997);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(989)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(989),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 990 transition  input  output  no-bypass 
    -- predecessors 653 
    -- successors 991 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4739_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_base_resize_ack_0, ack => cp_elements(990)); -- 
    sum_rename_req_4743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(990), ack => ptr_deref_1113_root_address_inst_req_0); -- 
    -- CP-element group 991 transition  input  output  no-bypass 
    -- predecessors 990 
    -- successors 992 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_root_address_inst_ack_0, ack => cp_elements(991)); -- 
    root_register_req_4748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(991), ack => ptr_deref_1113_addr_0_req_0); -- 
    -- CP-element group 992 fork  transition  input  no-bypass 
    -- predecessors 991 
    -- successors 988 993 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_word_addrgen/root_register_ack
      -- 
    root_register_ack_4749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_addr_0_ack_0, ack => cp_elements(992)); -- 
    -- CP-element group 993 transition  output  bypass 
    -- predecessors 992 
    -- successors 994 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/word_access/word_access_0/rr
      -- 
    cp_elements(993) <= cp_elements(992);
    rr_4759_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(993), ack => ptr_deref_1113_load_0_req_0); -- 
    -- CP-element group 994 transition  input  no-bypass 
    -- predecessors 993 
    -- successors 988 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_request/word_access/word_access_0/ra
      -- 
    ra_4760_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_0_ack_0, ack => cp_elements(994)); -- 
    -- CP-element group 995 transition  output  bypass 
    -- predecessors 988 
    -- successors 996 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/word_access/word_access_0/cr
      -- 
    cp_elements(995) <= cp_elements(988);
    cr_4770_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(995), ack => ptr_deref_1113_load_0_req_1); -- 
    -- CP-element group 996 transition  input  output  no-bypass 
    -- predecessors 995 
    -- successors 997 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/merge_req
      -- 
    ca_4771_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_0_ack_1, ack => cp_elements(996)); -- 
    merge_req_4772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(996), ack => ptr_deref_1113_gather_scatter_req_0); -- 
    -- CP-element group 997 transition  input  no-bypass 
    -- predecessors 996 
    -- successors 989 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1113_complete/merge_ack
      -- 
    merge_ack_4773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_gather_scatter_ack_0, ack => cp_elements(997)); -- 
    -- CP-element group 998 join  fork  transition  bypass 
    -- predecessors 1002 1004 
    -- successors 999 1005 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_active_
      -- 
    cpelement_group_998 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1002);
      predecessors(1) <= cp_elements(1004);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(998)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(998),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 999 join  fork  transition  bypass 
    -- predecessors 998 1007 
    -- successors 1061 1481 1781 2081 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1118_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1118_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1118_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_completed_
      -- 
    cpelement_group_999 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(998);
      predecessors(1) <= cp_elements(1007);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(999)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(999),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1000 transition  input  output  no-bypass 
    -- predecessors 732 
    -- successors 1001 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_base_resize_ack_0, ack => cp_elements(1000)); -- 
    sum_rename_req_4795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1000), ack => ptr_deref_1117_root_address_inst_req_0); -- 
    -- CP-element group 1001 transition  input  output  no-bypass 
    -- predecessors 1000 
    -- successors 1002 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_root_address_inst_ack_0, ack => cp_elements(1001)); -- 
    root_register_req_4800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1001), ack => ptr_deref_1117_addr_0_req_0); -- 
    -- CP-element group 1002 fork  transition  input  no-bypass 
    -- predecessors 1001 
    -- successors 998 1003 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_word_addrgen/root_register_ack
      -- 
    root_register_ack_4801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_addr_0_ack_0, ack => cp_elements(1002)); -- 
    -- CP-element group 1003 transition  output  bypass 
    -- predecessors 1002 
    -- successors 1004 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/word_access/word_access_0/rr
      -- 
    cp_elements(1003) <= cp_elements(1002);
    rr_4811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1003), ack => ptr_deref_1117_load_0_req_0); -- 
    -- CP-element group 1004 transition  input  no-bypass 
    -- predecessors 1003 
    -- successors 998 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_request/word_access/word_access_0/ra
      -- 
    ra_4812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_load_0_ack_0, ack => cp_elements(1004)); -- 
    -- CP-element group 1005 transition  output  bypass 
    -- predecessors 998 
    -- successors 1006 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1005) <= cp_elements(998);
    cr_4822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1005), ack => ptr_deref_1117_load_0_req_1); -- 
    -- CP-element group 1006 transition  input  output  no-bypass 
    -- predecessors 1005 
    -- successors 1007 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/merge_req
      -- 
    ca_4823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_load_0_ack_1, ack => cp_elements(1006)); -- 
    merge_req_4824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1006), ack => ptr_deref_1117_gather_scatter_req_0); -- 
    -- CP-element group 1007 transition  input  no-bypass 
    -- predecessors 1006 
    -- successors 999 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1117_complete/merge_ack
      -- 
    merge_ack_4825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1117_gather_scatter_ack_0, ack => cp_elements(1007)); -- 
    -- CP-element group 1008 join  fork  transition  bypass 
    -- predecessors 1012 1014 
    -- successors 1009 1015 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_active_
      -- 
    cpelement_group_1008 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1012);
      predecessors(1) <= cp_elements(1014);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1008)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1008),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1009 join  fork  transition  bypass 
    -- predecessors 1008 1017 
    -- successors 1076 1181 1286 1391 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1122_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1122_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1122_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_completed_
      -- 
    cpelement_group_1009 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1008);
      predecessors(1) <= cp_elements(1017);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1009)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1009),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1010 transition  input  output  no-bypass 
    -- predecessors 425 
    -- successors 1011 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4843_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_base_resize_ack_0, ack => cp_elements(1010)); -- 
    sum_rename_req_4847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1010), ack => ptr_deref_1121_root_address_inst_req_0); -- 
    -- CP-element group 1011 transition  input  output  no-bypass 
    -- predecessors 1010 
    -- successors 1012 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_root_address_inst_ack_0, ack => cp_elements(1011)); -- 
    root_register_req_4852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1011), ack => ptr_deref_1121_addr_0_req_0); -- 
    -- CP-element group 1012 fork  transition  input  no-bypass 
    -- predecessors 1011 
    -- successors 1008 1013 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_word_addrgen/root_register_ack
      -- 
    root_register_ack_4853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_addr_0_ack_0, ack => cp_elements(1012)); -- 
    -- CP-element group 1013 transition  output  bypass 
    -- predecessors 1012 
    -- successors 1014 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/word_access/word_access_0/rr
      -- 
    cp_elements(1013) <= cp_elements(1012);
    rr_4863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1013), ack => ptr_deref_1121_load_0_req_0); -- 
    -- CP-element group 1014 transition  input  no-bypass 
    -- predecessors 1013 
    -- successors 1008 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_request/word_access/word_access_0/ra
      -- 
    ra_4864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_load_0_ack_0, ack => cp_elements(1014)); -- 
    -- CP-element group 1015 transition  output  bypass 
    -- predecessors 1008 
    -- successors 1016 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1015) <= cp_elements(1008);
    cr_4874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1015), ack => ptr_deref_1121_load_0_req_1); -- 
    -- CP-element group 1016 transition  input  output  no-bypass 
    -- predecessors 1015 
    -- successors 1017 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/merge_req
      -- 
    ca_4875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_load_0_ack_1, ack => cp_elements(1016)); -- 
    merge_req_4876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1016), ack => ptr_deref_1121_gather_scatter_req_0); -- 
    -- CP-element group 1017 transition  input  no-bypass 
    -- predecessors 1016 
    -- successors 1009 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1121_complete/merge_ack
      -- 
    merge_ack_4877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1121_gather_scatter_ack_0, ack => cp_elements(1017)); -- 
    -- CP-element group 1018 join  fork  transition  bypass 
    -- predecessors 1022 1024 
    -- successors 1019 1025 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_active_
      -- 
    cpelement_group_1018 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1022);
      predecessors(1) <= cp_elements(1024);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1018)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1018),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1019 join  fork  transition  bypass 
    -- predecessors 1018 1027 
    -- successors 1077 1497 1797 2097 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1126_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1126_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1126_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_completed_
      -- 
    cpelement_group_1019 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1018);
      predecessors(1) <= cp_elements(1027);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1019)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1019),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1020 transition  input  output  no-bypass 
    -- predecessors 708 
    -- successors 1021 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_base_resize_ack_0, ack => cp_elements(1020)); -- 
    sum_rename_req_4899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1020), ack => ptr_deref_1125_root_address_inst_req_0); -- 
    -- CP-element group 1021 transition  input  output  no-bypass 
    -- predecessors 1020 
    -- successors 1022 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_word_addrgen/root_register_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_root_address_inst_ack_0, ack => cp_elements(1021)); -- 
    root_register_req_4904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1021), ack => ptr_deref_1125_addr_0_req_0); -- 
    -- CP-element group 1022 fork  transition  input  no-bypass 
    -- predecessors 1021 
    -- successors 1018 1023 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_word_addrgen/root_register_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_word_address_calculated
      -- 
    root_register_ack_4905_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_addr_0_ack_0, ack => cp_elements(1022)); -- 
    -- CP-element group 1023 transition  output  bypass 
    -- predecessors 1022 
    -- successors 1024 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/word_access/word_access_0/rr
      -- 
    cp_elements(1023) <= cp_elements(1022);
    rr_4915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1023), ack => ptr_deref_1125_load_0_req_0); -- 
    -- CP-element group 1024 transition  input  no-bypass 
    -- predecessors 1023 
    -- successors 1018 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_request/word_access/word_access_0/ra
      -- 
    ra_4916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_load_0_ack_0, ack => cp_elements(1024)); -- 
    -- CP-element group 1025 transition  output  bypass 
    -- predecessors 1018 
    -- successors 1026 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1025) <= cp_elements(1018);
    cr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1025), ack => ptr_deref_1125_load_0_req_1); -- 
    -- CP-element group 1026 transition  input  output  no-bypass 
    -- predecessors 1025 
    -- successors 1027 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/merge_req
      -- 
    ca_4927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_load_0_ack_1, ack => cp_elements(1026)); -- 
    merge_req_4928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1026), ack => ptr_deref_1125_gather_scatter_req_0); -- 
    -- CP-element group 1027 transition  input  no-bypass 
    -- predecessors 1026 
    -- successors 1019 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1125_complete/merge_ack
      -- 
    merge_ack_4929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_gather_scatter_ack_0, ack => cp_elements(1027)); -- 
    -- CP-element group 1028 join  fork  transition  bypass 
    -- predecessors 1032 1034 
    -- successors 1029 1035 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_active_
      -- 
    cpelement_group_1028 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1032);
      predecessors(1) <= cp_elements(1034);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1028)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1028),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1029 join  fork  transition  bypass 
    -- predecessors 1028 1037 
    -- successors 1085 1190 1295 1400 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1130_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1130_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1130_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_completed_
      -- 
    cpelement_group_1029 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1028);
      predecessors(1) <= cp_elements(1037);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1029)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1029),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1030 transition  input  output  no-bypass 
    -- predecessors 401 
    -- successors 1031 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4947_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1129_base_resize_ack_0, ack => cp_elements(1030)); -- 
    sum_rename_req_4951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1030), ack => ptr_deref_1129_root_address_inst_req_0); -- 
    -- CP-element group 1031 transition  input  output  no-bypass 
    -- predecessors 1030 
    -- successors 1032 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1129_root_address_inst_ack_0, ack => cp_elements(1031)); -- 
    root_register_req_4956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1031), ack => ptr_deref_1129_addr_0_req_0); -- 
    -- CP-element group 1032 fork  transition  input  no-bypass 
    -- predecessors 1031 
    -- successors 1028 1033 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_word_addrgen/root_register_ack
      -- 
    root_register_ack_4957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1129_addr_0_ack_0, ack => cp_elements(1032)); -- 
    -- CP-element group 1033 transition  output  bypass 
    -- predecessors 1032 
    -- successors 1034 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/word_access/word_access_0/rr
      -- 
    cp_elements(1033) <= cp_elements(1032);
    rr_4967_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1033), ack => ptr_deref_1129_load_0_req_0); -- 
    -- CP-element group 1034 transition  input  no-bypass 
    -- predecessors 1033 
    -- successors 1028 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_request/word_access/word_access_0/ra
      -- 
    ra_4968_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1129_load_0_ack_0, ack => cp_elements(1034)); -- 
    -- CP-element group 1035 transition  output  bypass 
    -- predecessors 1028 
    -- successors 1036 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1035) <= cp_elements(1028);
    cr_4978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1035), ack => ptr_deref_1129_load_0_req_1); -- 
    -- CP-element group 1036 transition  input  output  no-bypass 
    -- predecessors 1035 
    -- successors 1037 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/merge_req
      -- 
    ca_4979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1129_load_0_ack_1, ack => cp_elements(1036)); -- 
    merge_req_4980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1036), ack => ptr_deref_1129_gather_scatter_req_0); -- 
    -- CP-element group 1037 transition  input  no-bypass 
    -- predecessors 1036 
    -- successors 1029 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1129_complete/merge_ack
      -- 
    merge_ack_4981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1129_gather_scatter_ack_0, ack => cp_elements(1037)); -- 
    -- CP-element group 1038 join  fork  transition  bypass 
    -- predecessors 1042 1044 
    -- successors 1039 1045 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_active_
      -- 
    cpelement_group_1038 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1042);
      predecessors(1) <= cp_elements(1044);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1038)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1038),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1039 join  fork  transition  bypass 
    -- predecessors 1038 1047 
    -- successors 1086 1506 1806 2106 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1134_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1134_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1134_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_completed_
      -- 
    cpelement_group_1039 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1038);
      predecessors(1) <= cp_elements(1047);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1039)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1039),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1040 transition  input  output  no-bypass 
    -- predecessors 684 
    -- successors 1041 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_address_resized
      -- 
    base_resize_ack_4999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_base_resize_ack_0, ack => cp_elements(1040)); -- 
    sum_rename_req_5003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1040), ack => ptr_deref_1133_root_address_inst_req_0); -- 
    -- CP-element group 1041 transition  input  output  no-bypass 
    -- predecessors 1040 
    -- successors 1042 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_word_addrgen/root_register_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_root_address_calculated
      -- 
    sum_rename_ack_5004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_root_address_inst_ack_0, ack => cp_elements(1041)); -- 
    root_register_req_5008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1041), ack => ptr_deref_1133_addr_0_req_0); -- 
    -- CP-element group 1042 fork  transition  input  no-bypass 
    -- predecessors 1041 
    -- successors 1038 1043 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_word_addrgen/root_register_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_word_address_calculated
      -- 
    root_register_ack_5009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_addr_0_ack_0, ack => cp_elements(1042)); -- 
    -- CP-element group 1043 transition  output  bypass 
    -- predecessors 1042 
    -- successors 1044 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/word_access/word_access_0/rr
      -- 
    cp_elements(1043) <= cp_elements(1042);
    rr_5019_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1043), ack => ptr_deref_1133_load_0_req_0); -- 
    -- CP-element group 1044 transition  input  no-bypass 
    -- predecessors 1043 
    -- successors 1038 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_request/word_access/word_access_0/ra
      -- 
    ra_5020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_load_0_ack_0, ack => cp_elements(1044)); -- 
    -- CP-element group 1045 transition  output  bypass 
    -- predecessors 1038 
    -- successors 1046 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1045) <= cp_elements(1038);
    cr_5030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1045), ack => ptr_deref_1133_load_0_req_1); -- 
    -- CP-element group 1046 transition  input  output  no-bypass 
    -- predecessors 1045 
    -- successors 1047 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/merge_req
      -- 
    ca_5031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_load_0_ack_1, ack => cp_elements(1046)); -- 
    merge_req_5032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1046), ack => ptr_deref_1133_gather_scatter_req_0); -- 
    -- CP-element group 1047 transition  input  no-bypass 
    -- predecessors 1046 
    -- successors 1039 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1133_complete/merge_ack
      -- 
    merge_ack_5033_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1133_gather_scatter_ack_0, ack => cp_elements(1047)); -- 
    -- CP-element group 1048 join  fork  transition  no-bypass 
    -- predecessors 1051 1052 
    -- successors 1049 1053 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_trigger_
      -- 
    cpelement_group_1048 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1051);
      predecessors(1) <= cp_elements(1052);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1048)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1048),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1049 join  fork  transition  no-bypass 
    -- predecessors 1048 1054 
    -- successors 1050 1055 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_active_
      -- 
    cpelement_group_1049 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1048);
      predecessors(1) <= cp_elements(1054);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1049)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1049),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1050 join  transition  bypass 
    -- predecessors 1049 1056 
    -- successors 1066 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1146_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1146_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1146_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1139_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1139_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1139_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_completed_
      -- 
    cpelement_group_1050 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1049);
      predecessors(1) <= cp_elements(1056);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1050)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1050),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1051 transition  bypass 
    -- predecessors 969 
    -- successors 1048 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1136_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1136_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1136_active_
      -- 
    cp_elements(1051) <= cp_elements(969);
    -- CP-element group 1052 transition  bypass 
    -- predecessors 979 
    -- successors 1048 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1137_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1137_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1137_completed_
      -- 
    cp_elements(1052) <= cp_elements(979);
    -- CP-element group 1053 transition  output  bypass 
    -- predecessors 1048 
    -- successors 1054 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Sample/rr
      -- 
    cp_elements(1053) <= cp_elements(1048);
    rr_5049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1053), ack => binary_1138_inst_req_0); -- 
    -- CP-element group 1054 transition  input  no-bypass 
    -- predecessors 1053 
    -- successors 1049 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Sample/$exit
      -- 
    ra_5050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1138_inst_ack_0, ack => cp_elements(1054)); -- 
    -- CP-element group 1055 transition  output  bypass 
    -- predecessors 1049 
    -- successors 1056 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Update/cr
      -- 
    cp_elements(1055) <= cp_elements(1049);
    cr_5054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1055), ack => binary_1138_inst_req_1); -- 
    -- CP-element group 1056 transition  input  no-bypass 
    -- predecessors 1055 
    -- successors 1050 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1138_complete_Update/ca
      -- 
    ca_5055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1138_inst_ack_1, ack => cp_elements(1056)); -- 
    -- CP-element group 1057 join  fork  transition  no-bypass 
    -- predecessors 1060 1061 
    -- successors 1058 1062 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_trigger_
      -- 
    cpelement_group_1057 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1060);
      predecessors(1) <= cp_elements(1061);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1057)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1057),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1058 join  fork  transition  no-bypass 
    -- predecessors 1057 1063 
    -- successors 1059 1064 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_active_
      -- 
    cpelement_group_1058 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1057);
      predecessors(1) <= cp_elements(1063);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1058)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1058),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1059 join  transition  bypass 
    -- predecessors 1058 1065 
    -- successors 1066 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1147_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1147_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1144_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1144_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1144_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1147_trigger_
      -- 
    cpelement_group_1059 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1058);
      predecessors(1) <= cp_elements(1065);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1059)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1059),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1060 transition  bypass 
    -- predecessors 989 
    -- successors 1057 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1141_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1141_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1141_completed_
      -- 
    cp_elements(1060) <= cp_elements(989);
    -- CP-element group 1061 transition  bypass 
    -- predecessors 999 
    -- successors 1057 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1142_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1142_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1142_completed_
      -- 
    cp_elements(1061) <= cp_elements(999);
    -- CP-element group 1062 transition  output  bypass 
    -- predecessors 1057 
    -- successors 1063 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Sample/rr
      -- 
    cp_elements(1062) <= cp_elements(1057);
    rr_5071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1062), ack => binary_1143_inst_req_0); -- 
    -- CP-element group 1063 transition  input  no-bypass 
    -- predecessors 1062 
    -- successors 1058 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Sample/ra
      -- 
    ra_5072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1143_inst_ack_0, ack => cp_elements(1063)); -- 
    -- CP-element group 1064 transition  output  bypass 
    -- predecessors 1058 
    -- successors 1065 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Update/$entry
      -- 
    cp_elements(1064) <= cp_elements(1058);
    cr_5076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1064), ack => binary_1143_inst_req_1); -- 
    -- CP-element group 1065 transition  input  no-bypass 
    -- predecessors 1064 
    -- successors 1059 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1143_complete_Update/$exit
      -- 
    ca_5077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1143_inst_ack_1, ack => cp_elements(1065)); -- 
    -- CP-element group 1066 join  fork  transition  bypass 
    -- predecessors 1050 1059 
    -- successors 1067 1069 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_trigger_
      -- 
    cpelement_group_1066 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1050);
      predecessors(1) <= cp_elements(1059);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1066)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1066),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1067 join  fork  transition  no-bypass 
    -- predecessors 1066 1070 
    -- successors 1068 1071 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_active_
      -- 
    cpelement_group_1067 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1066);
      predecessors(1) <= cp_elements(1070);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1067)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1067),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1068 join  transition  no-bypass 
    -- predecessors 1067 1072 
    -- successors 1098 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1149_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1149_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1149_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1166_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1166_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1166_completed_
      -- 
    cpelement_group_1068 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1067);
      predecessors(1) <= cp_elements(1072);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1068)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1068),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1069 transition  output  bypass 
    -- predecessors 1066 
    -- successors 1070 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Sample/$entry
      -- 
    cp_elements(1069) <= cp_elements(1066);
    rr_5093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1069), ack => binary_1148_inst_req_0); -- 
    -- CP-element group 1070 transition  input  no-bypass 
    -- predecessors 1069 
    -- successors 1067 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Sample/ra
      -- 
    ra_5094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1148_inst_ack_0, ack => cp_elements(1070)); -- 
    -- CP-element group 1071 transition  output  bypass 
    -- predecessors 1067 
    -- successors 1072 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Update/cr
      -- 
    cp_elements(1071) <= cp_elements(1067);
    cr_5098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1071), ack => binary_1148_inst_req_1); -- 
    -- CP-element group 1072 transition  input  no-bypass 
    -- predecessors 1071 
    -- successors 1068 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1148_complete_Update/ca
      -- 
    ca_5099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1148_inst_ack_1, ack => cp_elements(1072)); -- 
    -- CP-element group 1073 join  fork  transition  no-bypass 
    -- predecessors 1076 1077 
    -- successors 1074 1078 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_trigger_
      -- 
    cpelement_group_1073 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1076);
      predecessors(1) <= cp_elements(1077);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1073)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1073),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1074 join  fork  transition  no-bypass 
    -- predecessors 1073 1079 
    -- successors 1075 1080 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_active_
      -- 
    cpelement_group_1074 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1073);
      predecessors(1) <= cp_elements(1079);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1074)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1074),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1075 join  transition  bypass 
    -- predecessors 1074 1081 
    -- successors 1091 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1154_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1154_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1154_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1161_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1161_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1161_completed_
      -- 
    cpelement_group_1075 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1074);
      predecessors(1) <= cp_elements(1081);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1075)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1075),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1076 transition  bypass 
    -- predecessors 1009 
    -- successors 1073 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1151_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1151_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1151_active_
      -- 
    cp_elements(1076) <= cp_elements(1009);
    -- CP-element group 1077 transition  bypass 
    -- predecessors 1019 
    -- successors 1073 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1152_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1152_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1152_completed_
      -- 
    cp_elements(1077) <= cp_elements(1019);
    -- CP-element group 1078 transition  output  bypass 
    -- predecessors 1073 
    -- successors 1079 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Sample/rr
      -- 
    cp_elements(1078) <= cp_elements(1073);
    rr_5115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1078), ack => binary_1153_inst_req_0); -- 
    -- CP-element group 1079 transition  input  no-bypass 
    -- predecessors 1078 
    -- successors 1074 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Sample/$exit
      -- 
    ra_5116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1153_inst_ack_0, ack => cp_elements(1079)); -- 
    -- CP-element group 1080 transition  output  bypass 
    -- predecessors 1074 
    -- successors 1081 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Update/cr
      -- 
    cp_elements(1080) <= cp_elements(1074);
    cr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1080), ack => binary_1153_inst_req_1); -- 
    -- CP-element group 1081 transition  input  no-bypass 
    -- predecessors 1080 
    -- successors 1075 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1153_complete_Update/$exit
      -- 
    ca_5121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1153_inst_ack_1, ack => cp_elements(1081)); -- 
    -- CP-element group 1082 join  fork  transition  no-bypass 
    -- predecessors 1085 1086 
    -- successors 1083 1087 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_trigger_
      -- 
    cpelement_group_1082 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1085);
      predecessors(1) <= cp_elements(1086);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1082)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1082),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1083 join  fork  transition  no-bypass 
    -- predecessors 1082 1088 
    -- successors 1084 1089 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_active_
      -- 
    cpelement_group_1083 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1082);
      predecessors(1) <= cp_elements(1088);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1083)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1083),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1084 join  transition  bypass 
    -- predecessors 1083 1090 
    -- successors 1091 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1159_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1159_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1159_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1162_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1162_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1162_completed_
      -- 
    cpelement_group_1084 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1083);
      predecessors(1) <= cp_elements(1090);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1084)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1084),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1085 transition  bypass 
    -- predecessors 1029 
    -- successors 1082 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1156_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1156_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1156_active_
      -- 
    cp_elements(1085) <= cp_elements(1029);
    -- CP-element group 1086 transition  bypass 
    -- predecessors 1039 
    -- successors 1082 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1157_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1157_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1157_completed_
      -- 
    cp_elements(1086) <= cp_elements(1039);
    -- CP-element group 1087 transition  output  bypass 
    -- predecessors 1082 
    -- successors 1088 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Sample/$entry
      -- 
    cp_elements(1087) <= cp_elements(1082);
    rr_5137_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1087), ack => binary_1158_inst_req_0); -- 
    -- CP-element group 1088 transition  input  no-bypass 
    -- predecessors 1087 
    -- successors 1083 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Sample/ra
      -- 
    ra_5138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1158_inst_ack_0, ack => cp_elements(1088)); -- 
    -- CP-element group 1089 transition  output  bypass 
    -- predecessors 1083 
    -- successors 1090 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Update/cr
      -- 
    cp_elements(1089) <= cp_elements(1083);
    cr_5142_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1089), ack => binary_1158_inst_req_1); -- 
    -- CP-element group 1090 transition  input  no-bypass 
    -- predecessors 1089 
    -- successors 1084 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1158_complete_Update/ca
      -- 
    ca_5143_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1158_inst_ack_1, ack => cp_elements(1090)); -- 
    -- CP-element group 1091 join  fork  transition  bypass 
    -- predecessors 1075 1084 
    -- successors 1092 1094 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_trigger_
      -- 
    cpelement_group_1091 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1075);
      predecessors(1) <= cp_elements(1084);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1091)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1091),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1092 join  fork  transition  no-bypass 
    -- predecessors 1091 1095 
    -- successors 1093 1096 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_active_
      -- 
    cpelement_group_1092 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1091);
      predecessors(1) <= cp_elements(1095);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1092)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1092),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1093 join  transition  no-bypass 
    -- predecessors 1092 1097 
    -- successors 1098 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1164_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1164_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1164_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1167_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1167_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1167_completed_
      -- 
    cpelement_group_1093 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1092);
      predecessors(1) <= cp_elements(1097);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1093)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1093),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1094 transition  output  bypass 
    -- predecessors 1091 
    -- successors 1095 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Sample/rr
      -- 
    cp_elements(1094) <= cp_elements(1091);
    rr_5159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1094), ack => binary_1163_inst_req_0); -- 
    -- CP-element group 1095 transition  input  no-bypass 
    -- predecessors 1094 
    -- successors 1092 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Sample/ra
      -- 
    ra_5160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1163_inst_ack_0, ack => cp_elements(1095)); -- 
    -- CP-element group 1096 transition  output  bypass 
    -- predecessors 1092 
    -- successors 1097 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Update/cr
      -- 
    cp_elements(1096) <= cp_elements(1092);
    cr_5164_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1096), ack => binary_1163_inst_req_1); -- 
    -- CP-element group 1097 transition  input  no-bypass 
    -- predecessors 1096 
    -- successors 1093 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1163_complete_Update/ca
      -- 
    ca_5165_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1163_inst_ack_1, ack => cp_elements(1097)); -- 
    -- CP-element group 1098 join  fork  transition  bypass 
    -- predecessors 1068 1093 
    -- successors 1099 1101 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_trigger_
      -- 
    cpelement_group_1098 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1068);
      predecessors(1) <= cp_elements(1093);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1098)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1098),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1099 join  fork  transition  no-bypass 
    -- predecessors 1098 1102 
    -- successors 1100 1103 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_active_
      -- 
    cpelement_group_1099 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1098);
      predecessors(1) <= cp_elements(1102);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1099)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1099),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1100 join  transition  no-bypass 
    -- predecessors 1099 1104 
    -- successors 1105 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1169_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1169_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1169_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1172_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1172_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1172_completed_
      -- 
    cpelement_group_1100 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1099);
      predecessors(1) <= cp_elements(1104);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1100)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1101 transition  output  bypass 
    -- predecessors 1098 
    -- successors 1102 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Sample/rr
      -- 
    cp_elements(1101) <= cp_elements(1098);
    rr_5181_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1101), ack => binary_1168_inst_req_0); -- 
    -- CP-element group 1102 transition  input  no-bypass 
    -- predecessors 1101 
    -- successors 1099 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Sample/ra
      -- 
    ra_5182_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1168_inst_ack_0, ack => cp_elements(1102)); -- 
    -- CP-element group 1103 transition  output  bypass 
    -- predecessors 1099 
    -- successors 1104 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Update/cr
      -- 
    cp_elements(1103) <= cp_elements(1099);
    cr_5186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1103), ack => binary_1168_inst_req_1); -- 
    -- CP-element group 1104 transition  input  no-bypass 
    -- predecessors 1103 
    -- successors 1100 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1168_complete_Update/ca
      -- 
    ca_5187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1168_inst_ack_1, ack => cp_elements(1104)); -- 
    -- CP-element group 1105 join  fork  transition  no-bypass 
    -- predecessors 1100 1108 
    -- successors 1106 1109 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_trigger_
      -- 
    cpelement_group_1105 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1100);
      predecessors(1) <= cp_elements(1108);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1105)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1105),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1106 join  fork  transition  bypass 
    -- predecessors 1105 1110 
    -- successors 1107 1111 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_active_
      -- 
    cpelement_group_1106 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1105);
      predecessors(1) <= cp_elements(1110);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1106)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1106),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1107 join  transition  bypass 
    -- predecessors 1106 1112 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1174_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1174_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1174_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_completed_
      -- 
    cpelement_group_1107 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1106);
      predecessors(1) <= cp_elements(1112);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1107)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1107),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1108 transition  bypass 
    -- predecessors 367 
    -- successors 1105 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1171_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1171_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1171_completed_
      -- 
    cp_elements(1108) <= cp_elements(367);
    -- CP-element group 1109 transition  output  bypass 
    -- predecessors 1105 
    -- successors 1110 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Sample/rr
      -- 
    cp_elements(1109) <= cp_elements(1105);
    rr_5203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1109), ack => binary_1173_inst_req_0); -- 
    -- CP-element group 1110 transition  input  no-bypass 
    -- predecessors 1109 
    -- successors 1106 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Sample/ra
      -- 
    ra_5204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1173_inst_ack_0, ack => cp_elements(1110)); -- 
    -- CP-element group 1111 transition  output  bypass 
    -- predecessors 1106 
    -- successors 1112 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Update/cr
      -- 
    cp_elements(1111) <= cp_elements(1106);
    cr_5208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1111), ack => binary_1173_inst_req_1); -- 
    -- CP-element group 1112 transition  input  no-bypass 
    -- predecessors 1111 
    -- successors 1107 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1173_complete_Update/ca
      -- 
    ca_5209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1173_inst_ack_1, ack => cp_elements(1112)); -- 
    -- CP-element group 1113 join  fork  transition  bypass 
    -- predecessors 1117 1119 
    -- successors 1114 1120 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_active_
      -- 
    cpelement_group_1113 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1117);
      predecessors(1) <= cp_elements(1119);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1113)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1114 join  fork  transition  bypass 
    -- predecessors 1113 1122 
    -- successors 1157 1537 1837 2137 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1178_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1178_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1178_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_completed_
      -- 
    cpelement_group_1114 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1113);
      predecessors(1) <= cp_elements(1122);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1114)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1114),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1115 transition  input  output  no-bypass 
    -- predecessors 817 
    -- successors 1116 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1177_base_resize_ack_0, ack => cp_elements(1115)); -- 
    sum_rename_req_5231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1115), ack => ptr_deref_1177_root_address_inst_req_0); -- 
    -- CP-element group 1116 transition  input  output  no-bypass 
    -- predecessors 1115 
    -- successors 1117 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1177_root_address_inst_ack_0, ack => cp_elements(1116)); -- 
    root_register_req_5236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1116), ack => ptr_deref_1177_addr_0_req_0); -- 
    -- CP-element group 1117 fork  transition  input  no-bypass 
    -- predecessors 1116 
    -- successors 1113 1118 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_word_addrgen/root_register_ack
      -- 
    root_register_ack_5237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1177_addr_0_ack_0, ack => cp_elements(1117)); -- 
    -- CP-element group 1118 transition  output  bypass 
    -- predecessors 1117 
    -- successors 1119 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/word_access/word_access_0/rr
      -- 
    cp_elements(1118) <= cp_elements(1117);
    rr_5247_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1118), ack => ptr_deref_1177_load_0_req_0); -- 
    -- CP-element group 1119 transition  input  no-bypass 
    -- predecessors 1118 
    -- successors 1113 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_request/word_access/word_access_0/ra
      -- 
    ra_5248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1177_load_0_ack_0, ack => cp_elements(1119)); -- 
    -- CP-element group 1120 transition  output  bypass 
    -- predecessors 1113 
    -- successors 1121 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1120) <= cp_elements(1113);
    cr_5258_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1120), ack => ptr_deref_1177_load_0_req_1); -- 
    -- CP-element group 1121 transition  input  output  no-bypass 
    -- predecessors 1120 
    -- successors 1122 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/merge_req
      -- 
    ca_5259_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1177_load_0_ack_1, ack => cp_elements(1121)); -- 
    merge_req_5260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1121), ack => ptr_deref_1177_gather_scatter_req_0); -- 
    -- CP-element group 1122 transition  input  no-bypass 
    -- predecessors 1121 
    -- successors 1114 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1177_complete/merge_ack
      -- 
    merge_ack_5261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1177_gather_scatter_ack_0, ack => cp_elements(1122)); -- 
    -- CP-element group 1123 join  fork  transition  bypass 
    -- predecessors 1127 1129 
    -- successors 1124 1130 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_active_
      -- 
    cpelement_group_1123 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1127);
      predecessors(1) <= cp_elements(1129);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1123)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1123),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1124 join  fork  transition  bypass 
    -- predecessors 1123 1132 
    -- successors 1166 1546 1846 2146 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1182_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1182_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1182_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_completed_
      -- 
    cpelement_group_1124 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1123);
      predecessors(1) <= cp_elements(1132);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1124)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1124),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1125 transition  input  output  no-bypass 
    -- predecessors 800 
    -- successors 1126 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5279_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_base_resize_ack_0, ack => cp_elements(1125)); -- 
    sum_rename_req_5283_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1125), ack => ptr_deref_1181_root_address_inst_req_0); -- 
    -- CP-element group 1126 transition  input  output  no-bypass 
    -- predecessors 1125 
    -- successors 1127 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5284_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_root_address_inst_ack_0, ack => cp_elements(1126)); -- 
    root_register_req_5288_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1126), ack => ptr_deref_1181_addr_0_req_0); -- 
    -- CP-element group 1127 fork  transition  input  no-bypass 
    -- predecessors 1126 
    -- successors 1123 1128 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_word_addrgen/root_register_ack
      -- 
    root_register_ack_5289_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_addr_0_ack_0, ack => cp_elements(1127)); -- 
    -- CP-element group 1128 transition  output  bypass 
    -- predecessors 1127 
    -- successors 1129 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/word_access/word_access_0/rr
      -- 
    cp_elements(1128) <= cp_elements(1127);
    rr_5299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1128), ack => ptr_deref_1181_load_0_req_0); -- 
    -- CP-element group 1129 transition  input  no-bypass 
    -- predecessors 1128 
    -- successors 1123 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_request/word_access/word_access_0/ra
      -- 
    ra_5300_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_load_0_ack_0, ack => cp_elements(1129)); -- 
    -- CP-element group 1130 transition  output  bypass 
    -- predecessors 1123 
    -- successors 1131 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1130) <= cp_elements(1123);
    cr_5310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1130), ack => ptr_deref_1181_load_0_req_1); -- 
    -- CP-element group 1131 transition  input  output  no-bypass 
    -- predecessors 1130 
    -- successors 1132 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/merge_req
      -- 
    ca_5311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_load_0_ack_1, ack => cp_elements(1131)); -- 
    merge_req_5312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1131), ack => ptr_deref_1181_gather_scatter_req_0); -- 
    -- CP-element group 1132 transition  input  no-bypass 
    -- predecessors 1131 
    -- successors 1124 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1181_complete/merge_ack
      -- 
    merge_ack_5313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_gather_scatter_ack_0, ack => cp_elements(1132)); -- 
    -- CP-element group 1133 join  fork  transition  bypass 
    -- predecessors 1137 1139 
    -- successors 1134 1140 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_active_
      -- 
    cpelement_group_1133 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1137);
      predecessors(1) <= cp_elements(1139);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1133)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1133),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1134 join  fork  transition  bypass 
    -- predecessors 1133 1142 
    -- successors 1182 1562 1862 2162 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1186_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1186_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1186_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_completed_
      -- 
    cpelement_group_1134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1133);
      predecessors(1) <= cp_elements(1142);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1134)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1135 transition  input  output  no-bypass 
    -- predecessors 783 
    -- successors 1136 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_base_resize_ack_0, ack => cp_elements(1135)); -- 
    sum_rename_req_5335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1135), ack => ptr_deref_1185_root_address_inst_req_0); -- 
    -- CP-element group 1136 transition  input  output  no-bypass 
    -- predecessors 1135 
    -- successors 1137 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_root_address_inst_ack_0, ack => cp_elements(1136)); -- 
    root_register_req_5340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1136), ack => ptr_deref_1185_addr_0_req_0); -- 
    -- CP-element group 1137 fork  transition  input  no-bypass 
    -- predecessors 1136 
    -- successors 1133 1138 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_word_addrgen/root_register_ack
      -- 
    root_register_ack_5341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_addr_0_ack_0, ack => cp_elements(1137)); -- 
    -- CP-element group 1138 transition  output  bypass 
    -- predecessors 1137 
    -- successors 1139 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/word_access/word_access_0/rr
      -- 
    cp_elements(1138) <= cp_elements(1137);
    rr_5351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1138), ack => ptr_deref_1185_load_0_req_0); -- 
    -- CP-element group 1139 transition  input  no-bypass 
    -- predecessors 1138 
    -- successors 1133 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_request/word_access/word_access_0/ra
      -- 
    ra_5352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_load_0_ack_0, ack => cp_elements(1139)); -- 
    -- CP-element group 1140 transition  output  bypass 
    -- predecessors 1133 
    -- successors 1141 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1140) <= cp_elements(1133);
    cr_5362_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1140), ack => ptr_deref_1185_load_0_req_1); -- 
    -- CP-element group 1141 transition  input  output  no-bypass 
    -- predecessors 1140 
    -- successors 1142 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/merge_req
      -- 
    ca_5363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_load_0_ack_1, ack => cp_elements(1141)); -- 
    merge_req_5364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1141), ack => ptr_deref_1185_gather_scatter_req_0); -- 
    -- CP-element group 1142 transition  input  no-bypass 
    -- predecessors 1141 
    -- successors 1134 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1185_complete/merge_ack
      -- 
    merge_ack_5365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1185_gather_scatter_ack_0, ack => cp_elements(1142)); -- 
    -- CP-element group 1143 join  fork  transition  bypass 
    -- predecessors 1147 1149 
    -- successors 1144 1150 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_active_
      -- 
    cpelement_group_1143 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1147);
      predecessors(1) <= cp_elements(1149);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1143)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1143),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1144 join  fork  transition  bypass 
    -- predecessors 1143 1152 
    -- successors 1191 1571 1871 2171 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1190_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1190_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1190_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_completed_
      -- 
    cpelement_group_1144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1143);
      predecessors(1) <= cp_elements(1152);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1144)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1145 transition  input  output  no-bypass 
    -- predecessors 766 
    -- successors 1146 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1189_base_resize_ack_0, ack => cp_elements(1145)); -- 
    sum_rename_req_5387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1145), ack => ptr_deref_1189_root_address_inst_req_0); -- 
    -- CP-element group 1146 transition  input  output  no-bypass 
    -- predecessors 1145 
    -- successors 1147 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1189_root_address_inst_ack_0, ack => cp_elements(1146)); -- 
    root_register_req_5392_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1146), ack => ptr_deref_1189_addr_0_req_0); -- 
    -- CP-element group 1147 fork  transition  input  no-bypass 
    -- predecessors 1146 
    -- successors 1143 1148 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_word_addrgen/root_register_ack
      -- 
    root_register_ack_5393_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1189_addr_0_ack_0, ack => cp_elements(1147)); -- 
    -- CP-element group 1148 transition  output  bypass 
    -- predecessors 1147 
    -- successors 1149 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/word_access/word_access_0/rr
      -- 
    cp_elements(1148) <= cp_elements(1147);
    rr_5403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1148), ack => ptr_deref_1189_load_0_req_0); -- 
    -- CP-element group 1149 transition  input  no-bypass 
    -- predecessors 1148 
    -- successors 1143 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_request/word_access/word_access_0/ra
      -- 
    ra_5404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1189_load_0_ack_0, ack => cp_elements(1149)); -- 
    -- CP-element group 1150 transition  output  bypass 
    -- predecessors 1143 
    -- successors 1151 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1150) <= cp_elements(1143);
    cr_5414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1150), ack => ptr_deref_1189_load_0_req_1); -- 
    -- CP-element group 1151 transition  input  output  no-bypass 
    -- predecessors 1150 
    -- successors 1152 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/merge_req
      -- 
    ca_5415_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1189_load_0_ack_1, ack => cp_elements(1151)); -- 
    merge_req_5416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1151), ack => ptr_deref_1189_gather_scatter_req_0); -- 
    -- CP-element group 1152 transition  input  no-bypass 
    -- predecessors 1151 
    -- successors 1144 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1189_complete/merge_ack
      -- 
    merge_ack_5417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1189_gather_scatter_ack_0, ack => cp_elements(1152)); -- 
    -- CP-element group 1153 join  fork  transition  no-bypass 
    -- predecessors 1156 1157 
    -- successors 1154 1158 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_trigger_
      -- 
    cpelement_group_1153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1156);
      predecessors(1) <= cp_elements(1157);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1153)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1154 join  fork  transition  no-bypass 
    -- predecessors 1153 1159 
    -- successors 1155 1160 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_active_
      -- 
    cpelement_group_1154 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1153);
      predecessors(1) <= cp_elements(1159);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1154)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1154),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1155 join  transition  bypass 
    -- predecessors 1154 1161 
    -- successors 1171 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1195_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1195_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1195_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1202_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1202_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1202_completed_
      -- 
    cpelement_group_1155 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1154);
      predecessors(1) <= cp_elements(1161);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1155)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1156 transition  bypass 
    -- predecessors 969 
    -- successors 1153 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1192_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1192_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1192_completed_
      -- 
    cp_elements(1156) <= cp_elements(969);
    -- CP-element group 1157 transition  bypass 
    -- predecessors 1114 
    -- successors 1153 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1193_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1193_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1193_completed_
      -- 
    cp_elements(1157) <= cp_elements(1114);
    -- CP-element group 1158 transition  output  bypass 
    -- predecessors 1153 
    -- successors 1159 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Sample/rr
      -- 
    cp_elements(1158) <= cp_elements(1153);
    rr_5433_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1158), ack => binary_1194_inst_req_0); -- 
    -- CP-element group 1159 transition  input  no-bypass 
    -- predecessors 1158 
    -- successors 1154 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Sample/ra
      -- 
    ra_5434_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1194_inst_ack_0, ack => cp_elements(1159)); -- 
    -- CP-element group 1160 transition  output  bypass 
    -- predecessors 1154 
    -- successors 1161 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Update/cr
      -- 
    cp_elements(1160) <= cp_elements(1154);
    cr_5438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1160), ack => binary_1194_inst_req_1); -- 
    -- CP-element group 1161 transition  input  no-bypass 
    -- predecessors 1160 
    -- successors 1155 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1194_complete_Update/ca
      -- 
    ca_5439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1194_inst_ack_1, ack => cp_elements(1161)); -- 
    -- CP-element group 1162 join  fork  transition  no-bypass 
    -- predecessors 1165 1166 
    -- successors 1163 1167 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_trigger_
      -- 
    cpelement_group_1162 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1165);
      predecessors(1) <= cp_elements(1166);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1162)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1162),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1163 join  fork  transition  no-bypass 
    -- predecessors 1162 1168 
    -- successors 1164 1169 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_active_
      -- 
    cpelement_group_1163 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1162);
      predecessors(1) <= cp_elements(1168);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1163)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1163),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1164 join  transition  bypass 
    -- predecessors 1163 1170 
    -- successors 1171 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1200_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1200_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1200_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1203_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1203_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1203_completed_
      -- 
    cpelement_group_1164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1163);
      predecessors(1) <= cp_elements(1170);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1164)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1165 transition  bypass 
    -- predecessors 989 
    -- successors 1162 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1197_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1197_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1197_completed_
      -- 
    cp_elements(1165) <= cp_elements(989);
    -- CP-element group 1166 transition  bypass 
    -- predecessors 1124 
    -- successors 1162 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1198_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1198_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1198_completed_
      -- 
    cp_elements(1166) <= cp_elements(1124);
    -- CP-element group 1167 transition  output  bypass 
    -- predecessors 1162 
    -- successors 1168 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Sample/rr
      -- 
    cp_elements(1167) <= cp_elements(1162);
    rr_5455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1167), ack => binary_1199_inst_req_0); -- 
    -- CP-element group 1168 transition  input  no-bypass 
    -- predecessors 1167 
    -- successors 1163 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Sample/ra
      -- 
    ra_5456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1199_inst_ack_0, ack => cp_elements(1168)); -- 
    -- CP-element group 1169 transition  output  bypass 
    -- predecessors 1163 
    -- successors 1170 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Update/cr
      -- 
    cp_elements(1169) <= cp_elements(1163);
    cr_5460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1169), ack => binary_1199_inst_req_1); -- 
    -- CP-element group 1170 transition  input  no-bypass 
    -- predecessors 1169 
    -- successors 1164 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1199_complete_Update/ca
      -- 
    ca_5461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1199_inst_ack_1, ack => cp_elements(1170)); -- 
    -- CP-element group 1171 join  fork  transition  bypass 
    -- predecessors 1155 1164 
    -- successors 1172 1174 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_trigger_
      -- 
    cpelement_group_1171 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1155);
      predecessors(1) <= cp_elements(1164);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1171)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1171),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1172 join  fork  transition  no-bypass 
    -- predecessors 1171 1175 
    -- successors 1173 1176 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_active_
      -- 
    cpelement_group_1172 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1171);
      predecessors(1) <= cp_elements(1175);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1172)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1172),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1173 join  transition  no-bypass 
    -- predecessors 1172 1177 
    -- successors 1203 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1205_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1205_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1205_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1222_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1222_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1222_completed_
      -- 
    cpelement_group_1173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1172);
      predecessors(1) <= cp_elements(1177);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1173)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1174 transition  output  bypass 
    -- predecessors 1171 
    -- successors 1175 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Sample/rr
      -- 
    cp_elements(1174) <= cp_elements(1171);
    rr_5477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1174), ack => binary_1204_inst_req_0); -- 
    -- CP-element group 1175 transition  input  no-bypass 
    -- predecessors 1174 
    -- successors 1172 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Sample/ra
      -- 
    ra_5478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1204_inst_ack_0, ack => cp_elements(1175)); -- 
    -- CP-element group 1176 transition  output  bypass 
    -- predecessors 1172 
    -- successors 1177 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Update/cr
      -- 
    cp_elements(1176) <= cp_elements(1172);
    cr_5482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1176), ack => binary_1204_inst_req_1); -- 
    -- CP-element group 1177 transition  input  no-bypass 
    -- predecessors 1176 
    -- successors 1173 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1204_complete_Update/ca
      -- 
    ca_5483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1204_inst_ack_1, ack => cp_elements(1177)); -- 
    -- CP-element group 1178 join  fork  transition  no-bypass 
    -- predecessors 1181 1182 
    -- successors 1179 1183 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_trigger_
      -- 
    cpelement_group_1178 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1181);
      predecessors(1) <= cp_elements(1182);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1178)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1178),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1179 join  fork  transition  no-bypass 
    -- predecessors 1178 1184 
    -- successors 1180 1185 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_active_
      -- 
    cpelement_group_1179 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1178);
      predecessors(1) <= cp_elements(1184);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1179)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1179),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1180 join  transition  bypass 
    -- predecessors 1179 1186 
    -- successors 1196 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1210_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1210_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1210_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1217_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1217_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1217_completed_
      -- 
    cpelement_group_1180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1179);
      predecessors(1) <= cp_elements(1186);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1180)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1181 transition  bypass 
    -- predecessors 1009 
    -- successors 1178 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1207_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1207_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1207_completed_
      -- 
    cp_elements(1181) <= cp_elements(1009);
    -- CP-element group 1182 transition  bypass 
    -- predecessors 1134 
    -- successors 1178 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1208_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1208_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1208_completed_
      -- 
    cp_elements(1182) <= cp_elements(1134);
    -- CP-element group 1183 transition  output  bypass 
    -- predecessors 1178 
    -- successors 1184 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Sample/rr
      -- 
    cp_elements(1183) <= cp_elements(1178);
    rr_5499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1183), ack => binary_1209_inst_req_0); -- 
    -- CP-element group 1184 transition  input  no-bypass 
    -- predecessors 1183 
    -- successors 1179 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Sample/ra
      -- 
    ra_5500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1209_inst_ack_0, ack => cp_elements(1184)); -- 
    -- CP-element group 1185 transition  output  bypass 
    -- predecessors 1179 
    -- successors 1186 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Update/cr
      -- 
    cp_elements(1185) <= cp_elements(1179);
    cr_5504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1185), ack => binary_1209_inst_req_1); -- 
    -- CP-element group 1186 transition  input  no-bypass 
    -- predecessors 1185 
    -- successors 1180 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1209_complete_Update/ca
      -- 
    ca_5505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1209_inst_ack_1, ack => cp_elements(1186)); -- 
    -- CP-element group 1187 join  fork  transition  no-bypass 
    -- predecessors 1190 1191 
    -- successors 1188 1192 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_trigger_
      -- 
    cpelement_group_1187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1190);
      predecessors(1) <= cp_elements(1191);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1187)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1188 join  fork  transition  no-bypass 
    -- predecessors 1187 1193 
    -- successors 1189 1194 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_active_
      -- 
    cpelement_group_1188 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1187);
      predecessors(1) <= cp_elements(1193);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1188)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1188),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1189 join  transition  bypass 
    -- predecessors 1188 1195 
    -- successors 1196 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1215_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1215_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1215_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1218_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1218_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1218_completed_
      -- 
    cpelement_group_1189 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1188);
      predecessors(1) <= cp_elements(1195);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1189)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1189),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1190 transition  bypass 
    -- predecessors 1029 
    -- successors 1187 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1212_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1212_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1212_completed_
      -- 
    cp_elements(1190) <= cp_elements(1029);
    -- CP-element group 1191 transition  bypass 
    -- predecessors 1144 
    -- successors 1187 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1213_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1213_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1213_completed_
      -- 
    cp_elements(1191) <= cp_elements(1144);
    -- CP-element group 1192 transition  output  bypass 
    -- predecessors 1187 
    -- successors 1193 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Sample/rr
      -- 
    cp_elements(1192) <= cp_elements(1187);
    rr_5521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1192), ack => binary_1214_inst_req_0); -- 
    -- CP-element group 1193 transition  input  no-bypass 
    -- predecessors 1192 
    -- successors 1188 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Sample/ra
      -- 
    ra_5522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1214_inst_ack_0, ack => cp_elements(1193)); -- 
    -- CP-element group 1194 transition  output  bypass 
    -- predecessors 1188 
    -- successors 1195 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Update/cr
      -- 
    cp_elements(1194) <= cp_elements(1188);
    cr_5526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1194), ack => binary_1214_inst_req_1); -- 
    -- CP-element group 1195 transition  input  no-bypass 
    -- predecessors 1194 
    -- successors 1189 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1214_complete_Update/ca
      -- 
    ca_5527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1214_inst_ack_1, ack => cp_elements(1195)); -- 
    -- CP-element group 1196 join  fork  transition  bypass 
    -- predecessors 1180 1189 
    -- successors 1197 1199 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_trigger_
      -- 
    cpelement_group_1196 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1180);
      predecessors(1) <= cp_elements(1189);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1196)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1196),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1197 join  fork  transition  no-bypass 
    -- predecessors 1196 1200 
    -- successors 1198 1201 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_active_
      -- 
    cpelement_group_1197 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1196);
      predecessors(1) <= cp_elements(1200);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1197)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1197),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1198 join  transition  no-bypass 
    -- predecessors 1197 1202 
    -- successors 1203 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1220_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1220_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1220_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1223_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1223_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1223_completed_
      -- 
    cpelement_group_1198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1197);
      predecessors(1) <= cp_elements(1202);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1198)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1199 transition  output  bypass 
    -- predecessors 1196 
    -- successors 1200 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Sample/rr
      -- 
    cp_elements(1199) <= cp_elements(1196);
    rr_5543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1199), ack => binary_1219_inst_req_0); -- 
    -- CP-element group 1200 transition  input  no-bypass 
    -- predecessors 1199 
    -- successors 1197 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Sample/ra
      -- 
    ra_5544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1219_inst_ack_0, ack => cp_elements(1200)); -- 
    -- CP-element group 1201 transition  output  bypass 
    -- predecessors 1197 
    -- successors 1202 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Update/cr
      -- 
    cp_elements(1201) <= cp_elements(1197);
    cr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1201), ack => binary_1219_inst_req_1); -- 
    -- CP-element group 1202 transition  input  no-bypass 
    -- predecessors 1201 
    -- successors 1198 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1219_complete_Update/ca
      -- 
    ca_5549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1219_inst_ack_1, ack => cp_elements(1202)); -- 
    -- CP-element group 1203 join  fork  transition  bypass 
    -- predecessors 1173 1198 
    -- successors 1204 1206 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_trigger_
      -- 
    cpelement_group_1203 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1173);
      predecessors(1) <= cp_elements(1198);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1203)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1203),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1204 join  fork  transition  no-bypass 
    -- predecessors 1203 1207 
    -- successors 1205 1208 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_active_
      -- 
    cpelement_group_1204 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1203);
      predecessors(1) <= cp_elements(1207);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1204)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1205 join  transition  no-bypass 
    -- predecessors 1204 1209 
    -- successors 1210 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1225_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1225_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1225_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1228_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1228_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1228_completed_
      -- 
    cpelement_group_1205 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1204);
      predecessors(1) <= cp_elements(1209);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1205)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1205),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1206 transition  output  bypass 
    -- predecessors 1203 
    -- successors 1207 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Sample/rr
      -- 
    cp_elements(1206) <= cp_elements(1203);
    rr_5565_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1206), ack => binary_1224_inst_req_0); -- 
    -- CP-element group 1207 transition  input  no-bypass 
    -- predecessors 1206 
    -- successors 1204 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Sample/ra
      -- 
    ra_5566_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1224_inst_ack_0, ack => cp_elements(1207)); -- 
    -- CP-element group 1208 transition  output  bypass 
    -- predecessors 1204 
    -- successors 1209 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Update/cr
      -- 
    cp_elements(1208) <= cp_elements(1204);
    cr_5570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1208), ack => binary_1224_inst_req_1); -- 
    -- CP-element group 1209 transition  input  no-bypass 
    -- predecessors 1208 
    -- successors 1205 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1224_complete_Update/ca
      -- 
    ca_5571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1224_inst_ack_1, ack => cp_elements(1209)); -- 
    -- CP-element group 1210 join  fork  transition  no-bypass 
    -- predecessors 1205 1213 
    -- successors 1211 1214 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_trigger_
      -- 
    cpelement_group_1210 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1205);
      predecessors(1) <= cp_elements(1213);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1210)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1210),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1211 join  fork  transition  bypass 
    -- predecessors 1210 1215 
    -- successors 1212 1216 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_active_
      -- 
    cpelement_group_1211 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1210);
      predecessors(1) <= cp_elements(1215);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1211)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1211),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1212 join  transition  bypass 
    -- predecessors 1211 1217 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1230_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1230_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1230_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_completed_
      -- 
    cpelement_group_1212 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1211);
      predecessors(1) <= cp_elements(1217);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1212)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1212),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1213 transition  bypass 
    -- predecessors 367 
    -- successors 1210 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1227_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1227_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1227_completed_
      -- 
    cp_elements(1213) <= cp_elements(367);
    -- CP-element group 1214 transition  output  bypass 
    -- predecessors 1210 
    -- successors 1215 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Sample/rr
      -- 
    cp_elements(1214) <= cp_elements(1210);
    rr_5587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1214), ack => binary_1229_inst_req_0); -- 
    -- CP-element group 1215 transition  input  no-bypass 
    -- predecessors 1214 
    -- successors 1211 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Sample/ra
      -- 
    ra_5588_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1229_inst_ack_0, ack => cp_elements(1215)); -- 
    -- CP-element group 1216 transition  output  bypass 
    -- predecessors 1211 
    -- successors 1217 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Update/cr
      -- 
    cp_elements(1216) <= cp_elements(1211);
    cr_5592_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1216), ack => binary_1229_inst_req_1); -- 
    -- CP-element group 1217 transition  input  no-bypass 
    -- predecessors 1216 
    -- successors 1212 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1229_complete_Update/ca
      -- 
    ca_5593_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1229_inst_ack_1, ack => cp_elements(1217)); -- 
    -- CP-element group 1218 join  fork  transition  bypass 
    -- predecessors 1222 1224 
    -- successors 1219 1225 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_active_
      -- 
    cpelement_group_1218 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1222);
      predecessors(1) <= cp_elements(1224);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1218)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1218),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1219 join  fork  transition  bypass 
    -- predecessors 1218 1227 
    -- successors 1262 1602 1902 2202 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1234_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1234_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1234_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_completed_
      -- 
    cpelement_group_1219 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1218);
      predecessors(1) <= cp_elements(1227);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1219)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1219),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1220 transition  input  output  no-bypass 
    -- predecessors 885 
    -- successors 1221 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1233_base_resize_ack_0, ack => cp_elements(1220)); -- 
    sum_rename_req_5615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1220), ack => ptr_deref_1233_root_address_inst_req_0); -- 
    -- CP-element group 1221 transition  input  output  no-bypass 
    -- predecessors 1220 
    -- successors 1222 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5616_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1233_root_address_inst_ack_0, ack => cp_elements(1221)); -- 
    root_register_req_5620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1221), ack => ptr_deref_1233_addr_0_req_0); -- 
    -- CP-element group 1222 fork  transition  input  no-bypass 
    -- predecessors 1221 
    -- successors 1218 1223 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_word_addrgen/root_register_ack
      -- 
    root_register_ack_5621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1233_addr_0_ack_0, ack => cp_elements(1222)); -- 
    -- CP-element group 1223 transition  output  bypass 
    -- predecessors 1222 
    -- successors 1224 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/word_access/word_access_0/rr
      -- 
    cp_elements(1223) <= cp_elements(1222);
    rr_5631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1223), ack => ptr_deref_1233_load_0_req_0); -- 
    -- CP-element group 1224 transition  input  no-bypass 
    -- predecessors 1223 
    -- successors 1218 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_request/word_access/word_access_0/ra
      -- 
    ra_5632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1233_load_0_ack_0, ack => cp_elements(1224)); -- 
    -- CP-element group 1225 transition  output  bypass 
    -- predecessors 1218 
    -- successors 1226 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1225) <= cp_elements(1218);
    cr_5642_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1225), ack => ptr_deref_1233_load_0_req_1); -- 
    -- CP-element group 1226 transition  input  output  no-bypass 
    -- predecessors 1225 
    -- successors 1227 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/merge_req
      -- 
    ca_5643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1233_load_0_ack_1, ack => cp_elements(1226)); -- 
    merge_req_5644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1226), ack => ptr_deref_1233_gather_scatter_req_0); -- 
    -- CP-element group 1227 transition  input  no-bypass 
    -- predecessors 1226 
    -- successors 1219 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1233_complete/merge_ack
      -- 
    merge_ack_5645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1233_gather_scatter_ack_0, ack => cp_elements(1227)); -- 
    -- CP-element group 1228 join  fork  transition  bypass 
    -- predecessors 1232 1234 
    -- successors 1229 1235 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_active_
      -- 
    cpelement_group_1228 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1232);
      predecessors(1) <= cp_elements(1234);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1228)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1228),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1229 join  fork  transition  bypass 
    -- predecessors 1228 1237 
    -- successors 1271 1611 1911 2211 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1238_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1238_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1238_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_completed_
      -- 
    cpelement_group_1229 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1228);
      predecessors(1) <= cp_elements(1237);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1229)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1229),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1230 transition  input  output  no-bypass 
    -- predecessors 868 
    -- successors 1231 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5663_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1237_base_resize_ack_0, ack => cp_elements(1230)); -- 
    sum_rename_req_5667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1230), ack => ptr_deref_1237_root_address_inst_req_0); -- 
    -- CP-element group 1231 transition  input  output  no-bypass 
    -- predecessors 1230 
    -- successors 1232 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1237_root_address_inst_ack_0, ack => cp_elements(1231)); -- 
    root_register_req_5672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1231), ack => ptr_deref_1237_addr_0_req_0); -- 
    -- CP-element group 1232 fork  transition  input  no-bypass 
    -- predecessors 1231 
    -- successors 1228 1233 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_word_addrgen/root_register_ack
      -- 
    root_register_ack_5673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1237_addr_0_ack_0, ack => cp_elements(1232)); -- 
    -- CP-element group 1233 transition  output  bypass 
    -- predecessors 1232 
    -- successors 1234 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/word_access/word_access_0/rr
      -- 
    cp_elements(1233) <= cp_elements(1232);
    rr_5683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1233), ack => ptr_deref_1237_load_0_req_0); -- 
    -- CP-element group 1234 transition  input  no-bypass 
    -- predecessors 1233 
    -- successors 1228 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_request/word_access/word_access_0/ra
      -- 
    ra_5684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1237_load_0_ack_0, ack => cp_elements(1234)); -- 
    -- CP-element group 1235 transition  output  bypass 
    -- predecessors 1228 
    -- successors 1236 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1235) <= cp_elements(1228);
    cr_5694_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1235), ack => ptr_deref_1237_load_0_req_1); -- 
    -- CP-element group 1236 transition  input  output  no-bypass 
    -- predecessors 1235 
    -- successors 1237 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/merge_req
      -- 
    ca_5695_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1237_load_0_ack_1, ack => cp_elements(1236)); -- 
    merge_req_5696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1236), ack => ptr_deref_1237_gather_scatter_req_0); -- 
    -- CP-element group 1237 transition  input  no-bypass 
    -- predecessors 1236 
    -- successors 1229 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1237_complete/merge_ack
      -- 
    merge_ack_5697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1237_gather_scatter_ack_0, ack => cp_elements(1237)); -- 
    -- CP-element group 1238 join  fork  transition  bypass 
    -- predecessors 1242 1244 
    -- successors 1239 1245 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_active_
      -- 
    cpelement_group_1238 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1242);
      predecessors(1) <= cp_elements(1244);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1238)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1238),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1239 join  fork  transition  bypass 
    -- predecessors 1238 1247 
    -- successors 1287 1627 1927 2227 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1242_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1242_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1242_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_completed_
      -- 
    cpelement_group_1239 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1238);
      predecessors(1) <= cp_elements(1247);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1239)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1239),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1240 transition  input  output  no-bypass 
    -- predecessors 851 
    -- successors 1241 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1241_base_resize_ack_0, ack => cp_elements(1240)); -- 
    sum_rename_req_5719_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1240), ack => ptr_deref_1241_root_address_inst_req_0); -- 
    -- CP-element group 1241 transition  input  output  no-bypass 
    -- predecessors 1240 
    -- successors 1242 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5720_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1241_root_address_inst_ack_0, ack => cp_elements(1241)); -- 
    root_register_req_5724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1241), ack => ptr_deref_1241_addr_0_req_0); -- 
    -- CP-element group 1242 fork  transition  input  no-bypass 
    -- predecessors 1241 
    -- successors 1238 1243 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_word_addrgen/root_register_ack
      -- 
    root_register_ack_5725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1241_addr_0_ack_0, ack => cp_elements(1242)); -- 
    -- CP-element group 1243 transition  output  bypass 
    -- predecessors 1242 
    -- successors 1244 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/word_access/word_access_0/rr
      -- 
    cp_elements(1243) <= cp_elements(1242);
    rr_5735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1243), ack => ptr_deref_1241_load_0_req_0); -- 
    -- CP-element group 1244 transition  input  no-bypass 
    -- predecessors 1243 
    -- successors 1238 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_request/word_access/word_access_0/ra
      -- 
    ra_5736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1241_load_0_ack_0, ack => cp_elements(1244)); -- 
    -- CP-element group 1245 transition  output  bypass 
    -- predecessors 1238 
    -- successors 1246 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1245) <= cp_elements(1238);
    cr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1245), ack => ptr_deref_1241_load_0_req_1); -- 
    -- CP-element group 1246 transition  input  output  no-bypass 
    -- predecessors 1245 
    -- successors 1247 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/merge_req
      -- 
    ca_5747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1241_load_0_ack_1, ack => cp_elements(1246)); -- 
    merge_req_5748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1246), ack => ptr_deref_1241_gather_scatter_req_0); -- 
    -- CP-element group 1247 transition  input  no-bypass 
    -- predecessors 1246 
    -- successors 1239 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1241_complete/merge_ack
      -- 
    merge_ack_5749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1241_gather_scatter_ack_0, ack => cp_elements(1247)); -- 
    -- CP-element group 1248 join  fork  transition  bypass 
    -- predecessors 1252 1254 
    -- successors 1249 1255 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_active_
      -- 
    cpelement_group_1248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1252);
      predecessors(1) <= cp_elements(1254);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1248)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1249 join  fork  transition  bypass 
    -- predecessors 1248 1257 
    -- successors 1296 1636 1936 2236 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1246_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1246_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1246_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_completed_
      -- 
    cpelement_group_1249 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1248);
      predecessors(1) <= cp_elements(1257);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1249)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1249),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1250 transition  input  output  no-bypass 
    -- predecessors 834 
    -- successors 1251 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1245_base_resize_ack_0, ack => cp_elements(1250)); -- 
    sum_rename_req_5771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1250), ack => ptr_deref_1245_root_address_inst_req_0); -- 
    -- CP-element group 1251 transition  input  output  no-bypass 
    -- predecessors 1250 
    -- successors 1252 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1245_root_address_inst_ack_0, ack => cp_elements(1251)); -- 
    root_register_req_5776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1251), ack => ptr_deref_1245_addr_0_req_0); -- 
    -- CP-element group 1252 fork  transition  input  no-bypass 
    -- predecessors 1251 
    -- successors 1248 1253 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_word_addrgen/root_register_ack
      -- 
    root_register_ack_5777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1245_addr_0_ack_0, ack => cp_elements(1252)); -- 
    -- CP-element group 1253 transition  output  bypass 
    -- predecessors 1252 
    -- successors 1254 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/word_access/word_access_0/rr
      -- 
    cp_elements(1253) <= cp_elements(1252);
    rr_5787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1253), ack => ptr_deref_1245_load_0_req_0); -- 
    -- CP-element group 1254 transition  input  no-bypass 
    -- predecessors 1253 
    -- successors 1248 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_request/word_access/word_access_0/ra
      -- 
    ra_5788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1245_load_0_ack_0, ack => cp_elements(1254)); -- 
    -- CP-element group 1255 transition  output  bypass 
    -- predecessors 1248 
    -- successors 1256 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1255) <= cp_elements(1248);
    cr_5798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1255), ack => ptr_deref_1245_load_0_req_1); -- 
    -- CP-element group 1256 transition  input  output  no-bypass 
    -- predecessors 1255 
    -- successors 1257 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/merge_req
      -- 
    ca_5799_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1245_load_0_ack_1, ack => cp_elements(1256)); -- 
    merge_req_5800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1256), ack => ptr_deref_1245_gather_scatter_req_0); -- 
    -- CP-element group 1257 transition  input  no-bypass 
    -- predecessors 1256 
    -- successors 1249 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1245_complete/merge_ack
      -- 
    merge_ack_5801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1245_gather_scatter_ack_0, ack => cp_elements(1257)); -- 
    -- CP-element group 1258 join  fork  transition  no-bypass 
    -- predecessors 1261 1262 
    -- successors 1259 1263 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_trigger_
      -- 
    cpelement_group_1258 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1261);
      predecessors(1) <= cp_elements(1262);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1258)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1258),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1259 join  fork  transition  no-bypass 
    -- predecessors 1258 1264 
    -- successors 1260 1265 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_active_
      -- 
    cpelement_group_1259 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1258);
      predecessors(1) <= cp_elements(1264);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1259)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1259),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1260 join  transition  bypass 
    -- predecessors 1259 1266 
    -- successors 1276 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1251_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1251_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1251_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1258_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1258_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1258_completed_
      -- 
    cpelement_group_1260 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1259);
      predecessors(1) <= cp_elements(1266);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1260)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1260),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1261 transition  bypass 
    -- predecessors 969 
    -- successors 1258 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1248_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1248_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1248_completed_
      -- 
    cp_elements(1261) <= cp_elements(969);
    -- CP-element group 1262 transition  bypass 
    -- predecessors 1219 
    -- successors 1258 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1249_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1249_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1249_completed_
      -- 
    cp_elements(1262) <= cp_elements(1219);
    -- CP-element group 1263 transition  output  bypass 
    -- predecessors 1258 
    -- successors 1264 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Sample/rr
      -- 
    cp_elements(1263) <= cp_elements(1258);
    rr_5817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1263), ack => binary_1250_inst_req_0); -- 
    -- CP-element group 1264 transition  input  no-bypass 
    -- predecessors 1263 
    -- successors 1259 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Sample/ra
      -- 
    ra_5818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1250_inst_ack_0, ack => cp_elements(1264)); -- 
    -- CP-element group 1265 transition  output  bypass 
    -- predecessors 1259 
    -- successors 1266 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Update/cr
      -- 
    cp_elements(1265) <= cp_elements(1259);
    cr_5822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1265), ack => binary_1250_inst_req_1); -- 
    -- CP-element group 1266 transition  input  no-bypass 
    -- predecessors 1265 
    -- successors 1260 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1250_complete_Update/ca
      -- 
    ca_5823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1250_inst_ack_1, ack => cp_elements(1266)); -- 
    -- CP-element group 1267 join  fork  transition  no-bypass 
    -- predecessors 1270 1271 
    -- successors 1268 1272 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_trigger_
      -- 
    cpelement_group_1267 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1270);
      predecessors(1) <= cp_elements(1271);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1267)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1267),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1268 join  fork  transition  no-bypass 
    -- predecessors 1267 1273 
    -- successors 1269 1274 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_active_
      -- 
    cpelement_group_1268 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1267);
      predecessors(1) <= cp_elements(1273);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1268)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1268),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1269 join  transition  bypass 
    -- predecessors 1268 1275 
    -- successors 1276 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1256_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1256_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1256_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1259_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1259_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1259_completed_
      -- 
    cpelement_group_1269 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1268);
      predecessors(1) <= cp_elements(1275);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1269)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1269),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1270 transition  bypass 
    -- predecessors 989 
    -- successors 1267 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1253_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1253_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1253_completed_
      -- 
    cp_elements(1270) <= cp_elements(989);
    -- CP-element group 1271 transition  bypass 
    -- predecessors 1229 
    -- successors 1267 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1254_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1254_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1254_completed_
      -- 
    cp_elements(1271) <= cp_elements(1229);
    -- CP-element group 1272 transition  output  bypass 
    -- predecessors 1267 
    -- successors 1273 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Sample/rr
      -- 
    cp_elements(1272) <= cp_elements(1267);
    rr_5839_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1272), ack => binary_1255_inst_req_0); -- 
    -- CP-element group 1273 transition  input  no-bypass 
    -- predecessors 1272 
    -- successors 1268 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Sample/ra
      -- 
    ra_5840_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1255_inst_ack_0, ack => cp_elements(1273)); -- 
    -- CP-element group 1274 transition  output  bypass 
    -- predecessors 1268 
    -- successors 1275 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Update/cr
      -- 
    cp_elements(1274) <= cp_elements(1268);
    cr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1274), ack => binary_1255_inst_req_1); -- 
    -- CP-element group 1275 transition  input  no-bypass 
    -- predecessors 1274 
    -- successors 1269 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1255_complete_Update/ca
      -- 
    ca_5845_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1255_inst_ack_1, ack => cp_elements(1275)); -- 
    -- CP-element group 1276 join  fork  transition  bypass 
    -- predecessors 1260 1269 
    -- successors 1277 1279 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_trigger_
      -- 
    cpelement_group_1276 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1260);
      predecessors(1) <= cp_elements(1269);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1276)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1276),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1277 join  fork  transition  no-bypass 
    -- predecessors 1276 1280 
    -- successors 1278 1281 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_active_
      -- 
    cpelement_group_1277 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1276);
      predecessors(1) <= cp_elements(1280);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1277)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1278 join  transition  no-bypass 
    -- predecessors 1277 1282 
    -- successors 1308 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1278_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1278_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1278_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1261_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1261_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1261_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_completed_
      -- 
    cpelement_group_1278 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1277);
      predecessors(1) <= cp_elements(1282);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1278)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1278),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1279 transition  output  bypass 
    -- predecessors 1276 
    -- successors 1280 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Sample/rr
      -- 
    cp_elements(1279) <= cp_elements(1276);
    rr_5861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1279), ack => binary_1260_inst_req_0); -- 
    -- CP-element group 1280 transition  input  no-bypass 
    -- predecessors 1279 
    -- successors 1277 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Sample/ra
      -- 
    ra_5862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1260_inst_ack_0, ack => cp_elements(1280)); -- 
    -- CP-element group 1281 transition  output  bypass 
    -- predecessors 1277 
    -- successors 1282 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Update/cr
      -- 
    cp_elements(1281) <= cp_elements(1277);
    cr_5866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1281), ack => binary_1260_inst_req_1); -- 
    -- CP-element group 1282 transition  input  no-bypass 
    -- predecessors 1281 
    -- successors 1278 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1260_complete_Update/ca
      -- 
    ca_5867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1260_inst_ack_1, ack => cp_elements(1282)); -- 
    -- CP-element group 1283 join  fork  transition  no-bypass 
    -- predecessors 1286 1287 
    -- successors 1284 1288 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_trigger_
      -- 
    cpelement_group_1283 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1286);
      predecessors(1) <= cp_elements(1287);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1283)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1283),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1284 join  fork  transition  no-bypass 
    -- predecessors 1283 1289 
    -- successors 1285 1290 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_active_
      -- 
    cpelement_group_1284 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1283);
      predecessors(1) <= cp_elements(1289);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1284)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1284),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1285 join  transition  bypass 
    -- predecessors 1284 1291 
    -- successors 1301 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1273_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1273_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1273_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1266_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1266_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1266_completed_
      -- 
    cpelement_group_1285 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1284);
      predecessors(1) <= cp_elements(1291);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1285)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1285),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1286 transition  bypass 
    -- predecessors 1009 
    -- successors 1283 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1263_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1263_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1263_completed_
      -- 
    cp_elements(1286) <= cp_elements(1009);
    -- CP-element group 1287 transition  bypass 
    -- predecessors 1239 
    -- successors 1283 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1264_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1264_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1264_completed_
      -- 
    cp_elements(1287) <= cp_elements(1239);
    -- CP-element group 1288 transition  output  bypass 
    -- predecessors 1283 
    -- successors 1289 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Sample/rr
      -- 
    cp_elements(1288) <= cp_elements(1283);
    rr_5883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1288), ack => binary_1265_inst_req_0); -- 
    -- CP-element group 1289 transition  input  no-bypass 
    -- predecessors 1288 
    -- successors 1284 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Sample/ra
      -- 
    ra_5884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1265_inst_ack_0, ack => cp_elements(1289)); -- 
    -- CP-element group 1290 transition  output  bypass 
    -- predecessors 1284 
    -- successors 1291 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Update/cr
      -- 
    cp_elements(1290) <= cp_elements(1284);
    cr_5888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1290), ack => binary_1265_inst_req_1); -- 
    -- CP-element group 1291 transition  input  no-bypass 
    -- predecessors 1290 
    -- successors 1285 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1265_complete_Update/ca
      -- 
    ca_5889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1265_inst_ack_1, ack => cp_elements(1291)); -- 
    -- CP-element group 1292 join  fork  transition  no-bypass 
    -- predecessors 1295 1296 
    -- successors 1293 1297 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_trigger_
      -- 
    cpelement_group_1292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1295);
      predecessors(1) <= cp_elements(1296);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1292)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1293 join  fork  transition  no-bypass 
    -- predecessors 1292 1298 
    -- successors 1294 1299 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_active_
      -- 
    cpelement_group_1293 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1292);
      predecessors(1) <= cp_elements(1298);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1293)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1293),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1294 join  transition  bypass 
    -- predecessors 1293 1300 
    -- successors 1301 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1271_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1271_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1271_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1274_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1274_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1274_completed_
      -- 
    cpelement_group_1294 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1293);
      predecessors(1) <= cp_elements(1300);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1294)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1294),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1295 transition  bypass 
    -- predecessors 1029 
    -- successors 1292 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1268_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1268_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1268_completed_
      -- 
    cp_elements(1295) <= cp_elements(1029);
    -- CP-element group 1296 transition  bypass 
    -- predecessors 1249 
    -- successors 1292 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1269_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1269_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1269_completed_
      -- 
    cp_elements(1296) <= cp_elements(1249);
    -- CP-element group 1297 transition  output  bypass 
    -- predecessors 1292 
    -- successors 1298 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Sample/rr
      -- 
    cp_elements(1297) <= cp_elements(1292);
    rr_5905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1297), ack => binary_1270_inst_req_0); -- 
    -- CP-element group 1298 transition  input  no-bypass 
    -- predecessors 1297 
    -- successors 1293 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Sample/ra
      -- 
    ra_5906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1270_inst_ack_0, ack => cp_elements(1298)); -- 
    -- CP-element group 1299 transition  output  bypass 
    -- predecessors 1293 
    -- successors 1300 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Update/cr
      -- 
    cp_elements(1299) <= cp_elements(1293);
    cr_5910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1299), ack => binary_1270_inst_req_1); -- 
    -- CP-element group 1300 transition  input  no-bypass 
    -- predecessors 1299 
    -- successors 1294 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1270_complete_Update/ca
      -- 
    ca_5911_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1270_inst_ack_1, ack => cp_elements(1300)); -- 
    -- CP-element group 1301 join  fork  transition  bypass 
    -- predecessors 1285 1294 
    -- successors 1302 1304 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_trigger_
      -- 
    cpelement_group_1301 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1285);
      predecessors(1) <= cp_elements(1294);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1301)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1301),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1302 join  fork  transition  no-bypass 
    -- predecessors 1301 1305 
    -- successors 1303 1306 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_active_
      -- 
    cpelement_group_1302 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1301);
      predecessors(1) <= cp_elements(1305);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1302)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1302),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1303 join  transition  no-bypass 
    -- predecessors 1302 1307 
    -- successors 1308 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1276_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1276_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1276_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1279_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1279_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1279_completed_
      -- 
    cpelement_group_1303 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1302);
      predecessors(1) <= cp_elements(1307);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1303)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1303),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1304 transition  output  bypass 
    -- predecessors 1301 
    -- successors 1305 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Sample/rr
      -- 
    cp_elements(1304) <= cp_elements(1301);
    rr_5927_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1304), ack => binary_1275_inst_req_0); -- 
    -- CP-element group 1305 transition  input  no-bypass 
    -- predecessors 1304 
    -- successors 1302 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Sample/ra
      -- 
    ra_5928_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1275_inst_ack_0, ack => cp_elements(1305)); -- 
    -- CP-element group 1306 transition  output  bypass 
    -- predecessors 1302 
    -- successors 1307 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Update/cr
      -- 
    cp_elements(1306) <= cp_elements(1302);
    cr_5932_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1306), ack => binary_1275_inst_req_1); -- 
    -- CP-element group 1307 transition  input  no-bypass 
    -- predecessors 1306 
    -- successors 1303 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1275_complete_Update/ca
      -- 
    ca_5933_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1275_inst_ack_1, ack => cp_elements(1307)); -- 
    -- CP-element group 1308 join  fork  transition  bypass 
    -- predecessors 1278 1303 
    -- successors 1309 1311 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_trigger_
      -- 
    cpelement_group_1308 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1278);
      predecessors(1) <= cp_elements(1303);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1308)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1309 join  fork  transition  no-bypass 
    -- predecessors 1308 1312 
    -- successors 1310 1313 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_active_
      -- 
    cpelement_group_1309 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1308);
      predecessors(1) <= cp_elements(1312);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1309)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1309),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1310 join  transition  no-bypass 
    -- predecessors 1309 1314 
    -- successors 1315 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1281_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1281_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1284_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1284_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1281_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1284_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_completed_
      -- 
    cpelement_group_1310 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1309);
      predecessors(1) <= cp_elements(1314);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1310)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1310),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1311 transition  output  bypass 
    -- predecessors 1308 
    -- successors 1312 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Sample/$entry
      -- 
    cp_elements(1311) <= cp_elements(1308);
    rr_5949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1311), ack => binary_1280_inst_req_0); -- 
    -- CP-element group 1312 transition  input  no-bypass 
    -- predecessors 1311 
    -- successors 1309 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Sample/ra
      -- 
    ra_5950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1280_inst_ack_0, ack => cp_elements(1312)); -- 
    -- CP-element group 1313 transition  output  bypass 
    -- predecessors 1309 
    -- successors 1314 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Update/cr
      -- 
    cp_elements(1313) <= cp_elements(1309);
    cr_5954_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1313), ack => binary_1280_inst_req_1); -- 
    -- CP-element group 1314 transition  input  no-bypass 
    -- predecessors 1313 
    -- successors 1310 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1280_complete_Update/ca
      -- 
    ca_5955_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1280_inst_ack_1, ack => cp_elements(1314)); -- 
    -- CP-element group 1315 join  fork  transition  no-bypass 
    -- predecessors 1310 1318 
    -- successors 1316 1319 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_trigger_
      -- 
    cpelement_group_1315 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1310);
      predecessors(1) <= cp_elements(1318);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1315)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1315),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1316 join  fork  transition  bypass 
    -- predecessors 1315 1320 
    -- successors 1317 1321 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_active_
      -- 
    cpelement_group_1316 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1315);
      predecessors(1) <= cp_elements(1320);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1316)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1316),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1317 join  transition  bypass 
    -- predecessors 1316 1322 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1286_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1286_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1286_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_completed_
      -- 
    cpelement_group_1317 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1316);
      predecessors(1) <= cp_elements(1322);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1317)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1317),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1318 transition  bypass 
    -- predecessors 367 
    -- successors 1315 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1283_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1283_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1283_completed_
      -- 
    cp_elements(1318) <= cp_elements(367);
    -- CP-element group 1319 transition  output  bypass 
    -- predecessors 1315 
    -- successors 1320 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Sample/rr
      -- 
    cp_elements(1319) <= cp_elements(1315);
    rr_5971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1319), ack => binary_1285_inst_req_0); -- 
    -- CP-element group 1320 transition  input  no-bypass 
    -- predecessors 1319 
    -- successors 1316 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Sample/$exit
      -- 
    ra_5972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1285_inst_ack_0, ack => cp_elements(1320)); -- 
    -- CP-element group 1321 transition  output  bypass 
    -- predecessors 1316 
    -- successors 1322 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Update/cr
      -- 
    cp_elements(1321) <= cp_elements(1316);
    cr_5976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1321), ack => binary_1285_inst_req_1); -- 
    -- CP-element group 1322 transition  input  no-bypass 
    -- predecessors 1321 
    -- successors 1317 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1285_complete_Update/ca
      -- 
    ca_5977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1285_inst_ack_1, ack => cp_elements(1322)); -- 
    -- CP-element group 1323 join  fork  transition  bypass 
    -- predecessors 1327 1329 
    -- successors 1324 1330 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_active_
      -- 
    cpelement_group_1323 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1327);
      predecessors(1) <= cp_elements(1329);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1323)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1323),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1324 join  fork  transition  bypass 
    -- predecessors 1323 1332 
    -- successors 1367 1667 1967 2267 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1290_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1290_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1290_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_completed_
      -- 
    cpelement_group_1324 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1323);
      predecessors(1) <= cp_elements(1332);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1324)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1324),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1325 transition  input  output  no-bypass 
    -- predecessors 953 
    -- successors 1326 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_5995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_base_resize_ack_0, ack => cp_elements(1325)); -- 
    sum_rename_req_5999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1325), ack => ptr_deref_1289_root_address_inst_req_0); -- 
    -- CP-element group 1326 transition  input  output  no-bypass 
    -- predecessors 1325 
    -- successors 1327 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_word_addrgen/root_register_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_root_address_calculated
      -- 
    sum_rename_ack_6000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_root_address_inst_ack_0, ack => cp_elements(1326)); -- 
    root_register_req_6004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1326), ack => ptr_deref_1289_addr_0_req_0); -- 
    -- CP-element group 1327 fork  transition  input  no-bypass 
    -- predecessors 1326 
    -- successors 1323 1328 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_word_addrgen/root_register_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_word_addrgen/$exit
      -- 
    root_register_ack_6005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_addr_0_ack_0, ack => cp_elements(1327)); -- 
    -- CP-element group 1328 transition  output  bypass 
    -- predecessors 1327 
    -- successors 1329 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/word_access/word_access_0/$entry
      -- 
    cp_elements(1328) <= cp_elements(1327);
    rr_6015_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1328), ack => ptr_deref_1289_load_0_req_0); -- 
    -- CP-element group 1329 transition  input  no-bypass 
    -- predecessors 1328 
    -- successors 1323 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_request/word_access/word_access_0/ra
      -- 
    ra_6016_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_load_0_ack_0, ack => cp_elements(1329)); -- 
    -- CP-element group 1330 transition  output  bypass 
    -- predecessors 1323 
    -- successors 1331 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/$entry
      -- 
    cp_elements(1330) <= cp_elements(1323);
    cr_6026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1330), ack => ptr_deref_1289_load_0_req_1); -- 
    -- CP-element group 1331 transition  input  output  no-bypass 
    -- predecessors 1330 
    -- successors 1332 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/merge_req
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/word_access/word_access_0/$exit
      -- 
    ca_6027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_load_0_ack_1, ack => cp_elements(1331)); -- 
    merge_req_6028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1331), ack => ptr_deref_1289_gather_scatter_req_0); -- 
    -- CP-element group 1332 transition  input  no-bypass 
    -- predecessors 1331 
    -- successors 1324 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1289_complete/merge_ack
      -- 
    merge_ack_6029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_gather_scatter_ack_0, ack => cp_elements(1332)); -- 
    -- CP-element group 1333 join  fork  transition  bypass 
    -- predecessors 1337 1339 
    -- successors 1334 1340 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_active_
      -- 
    cpelement_group_1333 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1337);
      predecessors(1) <= cp_elements(1339);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1333)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1333),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1334 join  fork  transition  bypass 
    -- predecessors 1333 1342 
    -- successors 1376 1676 1976 2276 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1294_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1294_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1294_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_completed_
      -- 
    cpelement_group_1334 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1333);
      predecessors(1) <= cp_elements(1342);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1334)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1334),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1335 transition  input  output  no-bypass 
    -- predecessors 936 
    -- successors 1336 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6047_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1293_base_resize_ack_0, ack => cp_elements(1335)); -- 
    sum_rename_req_6051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1335), ack => ptr_deref_1293_root_address_inst_req_0); -- 
    -- CP-element group 1336 transition  input  output  no-bypass 
    -- predecessors 1335 
    -- successors 1337 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6052_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1293_root_address_inst_ack_0, ack => cp_elements(1336)); -- 
    root_register_req_6056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1336), ack => ptr_deref_1293_addr_0_req_0); -- 
    -- CP-element group 1337 fork  transition  input  no-bypass 
    -- predecessors 1336 
    -- successors 1333 1338 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_word_addrgen/root_register_ack
      -- 
    root_register_ack_6057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1293_addr_0_ack_0, ack => cp_elements(1337)); -- 
    -- CP-element group 1338 transition  output  bypass 
    -- predecessors 1337 
    -- successors 1339 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/word_access/word_access_0/rr
      -- 
    cp_elements(1338) <= cp_elements(1337);
    rr_6067_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1338), ack => ptr_deref_1293_load_0_req_0); -- 
    -- CP-element group 1339 transition  input  no-bypass 
    -- predecessors 1338 
    -- successors 1333 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_request/word_access/word_access_0/ra
      -- 
    ra_6068_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1293_load_0_ack_0, ack => cp_elements(1339)); -- 
    -- CP-element group 1340 transition  output  bypass 
    -- predecessors 1333 
    -- successors 1341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1340) <= cp_elements(1333);
    cr_6078_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1340), ack => ptr_deref_1293_load_0_req_1); -- 
    -- CP-element group 1341 transition  input  output  no-bypass 
    -- predecessors 1340 
    -- successors 1342 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/merge_req
      -- 
    ca_6079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1293_load_0_ack_1, ack => cp_elements(1341)); -- 
    merge_req_6080_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1341), ack => ptr_deref_1293_gather_scatter_req_0); -- 
    -- CP-element group 1342 transition  input  no-bypass 
    -- predecessors 1341 
    -- successors 1334 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1293_complete/merge_ack
      -- 
    merge_ack_6081_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1293_gather_scatter_ack_0, ack => cp_elements(1342)); -- 
    -- CP-element group 1343 join  fork  transition  bypass 
    -- predecessors 1347 1349 
    -- successors 1344 1350 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_active_
      -- 
    cpelement_group_1343 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1347);
      predecessors(1) <= cp_elements(1349);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1343)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1343),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1344 join  fork  transition  bypass 
    -- predecessors 1343 1352 
    -- successors 1392 1692 1992 2292 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1298_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1298_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1298_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_completed_
      -- 
    cpelement_group_1344 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1343);
      predecessors(1) <= cp_elements(1352);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1344)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1344),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1345 transition  input  output  no-bypass 
    -- predecessors 919 
    -- successors 1346 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1297_base_resize_ack_0, ack => cp_elements(1345)); -- 
    sum_rename_req_6103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1345), ack => ptr_deref_1297_root_address_inst_req_0); -- 
    -- CP-element group 1346 transition  input  output  no-bypass 
    -- predecessors 1345 
    -- successors 1347 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1297_root_address_inst_ack_0, ack => cp_elements(1346)); -- 
    root_register_req_6108_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1346), ack => ptr_deref_1297_addr_0_req_0); -- 
    -- CP-element group 1347 fork  transition  input  no-bypass 
    -- predecessors 1346 
    -- successors 1343 1348 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_word_addrgen/root_register_ack
      -- 
    root_register_ack_6109_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1297_addr_0_ack_0, ack => cp_elements(1347)); -- 
    -- CP-element group 1348 transition  output  bypass 
    -- predecessors 1347 
    -- successors 1349 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/word_access/word_access_0/rr
      -- 
    cp_elements(1348) <= cp_elements(1347);
    rr_6119_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1348), ack => ptr_deref_1297_load_0_req_0); -- 
    -- CP-element group 1349 transition  input  no-bypass 
    -- predecessors 1348 
    -- successors 1343 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_request/word_access/word_access_0/ra
      -- 
    ra_6120_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1297_load_0_ack_0, ack => cp_elements(1349)); -- 
    -- CP-element group 1350 transition  output  bypass 
    -- predecessors 1343 
    -- successors 1351 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1350) <= cp_elements(1343);
    cr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1350), ack => ptr_deref_1297_load_0_req_1); -- 
    -- CP-element group 1351 transition  input  output  no-bypass 
    -- predecessors 1350 
    -- successors 1352 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/merge_req
      -- 
    ca_6131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1297_load_0_ack_1, ack => cp_elements(1351)); -- 
    merge_req_6132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1351), ack => ptr_deref_1297_gather_scatter_req_0); -- 
    -- CP-element group 1352 transition  input  no-bypass 
    -- predecessors 1351 
    -- successors 1344 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1297_complete/merge_ack
      -- 
    merge_ack_6133_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1297_gather_scatter_ack_0, ack => cp_elements(1352)); -- 
    -- CP-element group 1353 join  fork  transition  bypass 
    -- predecessors 1357 1359 
    -- successors 1354 1360 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_active_
      -- 
    cpelement_group_1353 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1357);
      predecessors(1) <= cp_elements(1359);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1353)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1353),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1354 join  fork  transition  bypass 
    -- predecessors 1353 1362 
    -- successors 1401 1701 2001 2301 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1302_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1302_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1302_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_completed_
      -- 
    cpelement_group_1354 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1353);
      predecessors(1) <= cp_elements(1362);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1354)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1354),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1355 transition  input  output  no-bypass 
    -- predecessors 902 
    -- successors 1356 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1301_base_resize_ack_0, ack => cp_elements(1355)); -- 
    sum_rename_req_6155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1355), ack => ptr_deref_1301_root_address_inst_req_0); -- 
    -- CP-element group 1356 transition  input  output  no-bypass 
    -- predecessors 1355 
    -- successors 1357 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1301_root_address_inst_ack_0, ack => cp_elements(1356)); -- 
    root_register_req_6160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1356), ack => ptr_deref_1301_addr_0_req_0); -- 
    -- CP-element group 1357 fork  transition  input  no-bypass 
    -- predecessors 1356 
    -- successors 1353 1358 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_word_addrgen/root_register_ack
      -- 
    root_register_ack_6161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1301_addr_0_ack_0, ack => cp_elements(1357)); -- 
    -- CP-element group 1358 transition  output  bypass 
    -- predecessors 1357 
    -- successors 1359 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/word_access/word_access_0/rr
      -- 
    cp_elements(1358) <= cp_elements(1357);
    rr_6171_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1358), ack => ptr_deref_1301_load_0_req_0); -- 
    -- CP-element group 1359 transition  input  no-bypass 
    -- predecessors 1358 
    -- successors 1353 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_request/word_access/word_access_0/ra
      -- 
    ra_6172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1301_load_0_ack_0, ack => cp_elements(1359)); -- 
    -- CP-element group 1360 transition  output  bypass 
    -- predecessors 1353 
    -- successors 1361 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1360) <= cp_elements(1353);
    cr_6182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1360), ack => ptr_deref_1301_load_0_req_1); -- 
    -- CP-element group 1361 transition  input  output  no-bypass 
    -- predecessors 1360 
    -- successors 1362 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/merge_req
      -- 
    ca_6183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1301_load_0_ack_1, ack => cp_elements(1361)); -- 
    merge_req_6184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1361), ack => ptr_deref_1301_gather_scatter_req_0); -- 
    -- CP-element group 1362 transition  input  no-bypass 
    -- predecessors 1361 
    -- successors 1354 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1301_complete/merge_ack
      -- 
    merge_ack_6185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1301_gather_scatter_ack_0, ack => cp_elements(1362)); -- 
    -- CP-element group 1363 join  fork  transition  no-bypass 
    -- predecessors 1366 1367 
    -- successors 1364 1368 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_trigger_
      -- 
    cpelement_group_1363 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1366);
      predecessors(1) <= cp_elements(1367);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1363)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1363),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1364 join  fork  transition  no-bypass 
    -- predecessors 1363 1369 
    -- successors 1365 1370 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_active_
      -- 
    cpelement_group_1364 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1363);
      predecessors(1) <= cp_elements(1369);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1364)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1364),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1365 join  transition  bypass 
    -- predecessors 1364 1371 
    -- successors 1381 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1307_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1307_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1307_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1314_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1314_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1314_completed_
      -- 
    cpelement_group_1365 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1364);
      predecessors(1) <= cp_elements(1371);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1365)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1365),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1366 transition  bypass 
    -- predecessors 969 
    -- successors 1363 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1304_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1304_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1304_completed_
      -- 
    cp_elements(1366) <= cp_elements(969);
    -- CP-element group 1367 transition  bypass 
    -- predecessors 1324 
    -- successors 1363 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1305_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1305_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1305_completed_
      -- 
    cp_elements(1367) <= cp_elements(1324);
    -- CP-element group 1368 transition  output  bypass 
    -- predecessors 1363 
    -- successors 1369 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Sample/rr
      -- 
    cp_elements(1368) <= cp_elements(1363);
    rr_6201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1368), ack => binary_1306_inst_req_0); -- 
    -- CP-element group 1369 transition  input  no-bypass 
    -- predecessors 1368 
    -- successors 1364 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Sample/ra
      -- 
    ra_6202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1306_inst_ack_0, ack => cp_elements(1369)); -- 
    -- CP-element group 1370 transition  output  bypass 
    -- predecessors 1364 
    -- successors 1371 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Update/cr
      -- 
    cp_elements(1370) <= cp_elements(1364);
    cr_6206_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1370), ack => binary_1306_inst_req_1); -- 
    -- CP-element group 1371 transition  input  no-bypass 
    -- predecessors 1370 
    -- successors 1365 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1306_complete_Update/ca
      -- 
    ca_6207_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1306_inst_ack_1, ack => cp_elements(1371)); -- 
    -- CP-element group 1372 join  fork  transition  no-bypass 
    -- predecessors 1375 1376 
    -- successors 1373 1377 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_trigger_
      -- 
    cpelement_group_1372 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1375);
      predecessors(1) <= cp_elements(1376);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1372)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1372),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1373 join  fork  transition  no-bypass 
    -- predecessors 1372 1378 
    -- successors 1374 1379 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_active_
      -- 
    cpelement_group_1373 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1372);
      predecessors(1) <= cp_elements(1378);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1373)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1373),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1374 join  transition  bypass 
    -- predecessors 1373 1380 
    -- successors 1381 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1312_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1312_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1312_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1315_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1315_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1315_completed_
      -- 
    cpelement_group_1374 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1373);
      predecessors(1) <= cp_elements(1380);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1374)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1374),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1375 transition  bypass 
    -- predecessors 989 
    -- successors 1372 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1309_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1309_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1309_completed_
      -- 
    cp_elements(1375) <= cp_elements(989);
    -- CP-element group 1376 transition  bypass 
    -- predecessors 1334 
    -- successors 1372 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1310_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1310_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1310_completed_
      -- 
    cp_elements(1376) <= cp_elements(1334);
    -- CP-element group 1377 transition  output  bypass 
    -- predecessors 1372 
    -- successors 1378 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Sample/rr
      -- 
    cp_elements(1377) <= cp_elements(1372);
    rr_6223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1377), ack => binary_1311_inst_req_0); -- 
    -- CP-element group 1378 transition  input  no-bypass 
    -- predecessors 1377 
    -- successors 1373 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Sample/ra
      -- 
    ra_6224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1311_inst_ack_0, ack => cp_elements(1378)); -- 
    -- CP-element group 1379 transition  output  bypass 
    -- predecessors 1373 
    -- successors 1380 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Update/cr
      -- 
    cp_elements(1379) <= cp_elements(1373);
    cr_6228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1379), ack => binary_1311_inst_req_1); -- 
    -- CP-element group 1380 transition  input  no-bypass 
    -- predecessors 1379 
    -- successors 1374 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1311_complete_Update/ca
      -- 
    ca_6229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1311_inst_ack_1, ack => cp_elements(1380)); -- 
    -- CP-element group 1381 join  fork  transition  bypass 
    -- predecessors 1365 1374 
    -- successors 1382 1384 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_trigger_
      -- 
    cpelement_group_1381 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1365);
      predecessors(1) <= cp_elements(1374);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1381)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1381),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1382 join  fork  transition  no-bypass 
    -- predecessors 1381 1385 
    -- successors 1383 1386 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_active_
      -- 
    cpelement_group_1382 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1381);
      predecessors(1) <= cp_elements(1385);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1382)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1382),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1383 join  transition  no-bypass 
    -- predecessors 1382 1387 
    -- successors 1413 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1317_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1317_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1317_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1334_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1334_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1334_completed_
      -- 
    cpelement_group_1383 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1382);
      predecessors(1) <= cp_elements(1387);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1383)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1383),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1384 transition  output  bypass 
    -- predecessors 1381 
    -- successors 1385 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Sample/rr
      -- 
    cp_elements(1384) <= cp_elements(1381);
    rr_6245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1384), ack => binary_1316_inst_req_0); -- 
    -- CP-element group 1385 transition  input  no-bypass 
    -- predecessors 1384 
    -- successors 1382 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Sample/ra
      -- 
    ra_6246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1316_inst_ack_0, ack => cp_elements(1385)); -- 
    -- CP-element group 1386 transition  output  bypass 
    -- predecessors 1382 
    -- successors 1387 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Update/cr
      -- 
    cp_elements(1386) <= cp_elements(1382);
    cr_6250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1386), ack => binary_1316_inst_req_1); -- 
    -- CP-element group 1387 transition  input  no-bypass 
    -- predecessors 1386 
    -- successors 1383 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1316_complete_Update/ca
      -- 
    ca_6251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1316_inst_ack_1, ack => cp_elements(1387)); -- 
    -- CP-element group 1388 join  fork  transition  no-bypass 
    -- predecessors 1391 1392 
    -- successors 1389 1393 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_trigger_
      -- 
    cpelement_group_1388 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1391);
      predecessors(1) <= cp_elements(1392);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1388)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1388),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1389 join  fork  transition  no-bypass 
    -- predecessors 1388 1394 
    -- successors 1390 1395 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_active_
      -- 
    cpelement_group_1389 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1388);
      predecessors(1) <= cp_elements(1394);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1389)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1389),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1390 join  transition  bypass 
    -- predecessors 1389 1396 
    -- successors 1406 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1322_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1322_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1322_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1329_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1329_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1329_completed_
      -- 
    cpelement_group_1390 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1389);
      predecessors(1) <= cp_elements(1396);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1390)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1390),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1391 transition  bypass 
    -- predecessors 1009 
    -- successors 1388 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1319_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1319_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1319_completed_
      -- 
    cp_elements(1391) <= cp_elements(1009);
    -- CP-element group 1392 transition  bypass 
    -- predecessors 1344 
    -- successors 1388 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1320_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1320_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1320_completed_
      -- 
    cp_elements(1392) <= cp_elements(1344);
    -- CP-element group 1393 transition  output  bypass 
    -- predecessors 1388 
    -- successors 1394 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Sample/rr
      -- 
    cp_elements(1393) <= cp_elements(1388);
    rr_6267_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1393), ack => binary_1321_inst_req_0); -- 
    -- CP-element group 1394 transition  input  no-bypass 
    -- predecessors 1393 
    -- successors 1389 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Sample/ra
      -- 
    ra_6268_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1321_inst_ack_0, ack => cp_elements(1394)); -- 
    -- CP-element group 1395 transition  output  bypass 
    -- predecessors 1389 
    -- successors 1396 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Update/cr
      -- 
    cp_elements(1395) <= cp_elements(1389);
    cr_6272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1395), ack => binary_1321_inst_req_1); -- 
    -- CP-element group 1396 transition  input  no-bypass 
    -- predecessors 1395 
    -- successors 1390 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1321_complete_Update/ca
      -- 
    ca_6273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1321_inst_ack_1, ack => cp_elements(1396)); -- 
    -- CP-element group 1397 join  fork  transition  no-bypass 
    -- predecessors 1400 1401 
    -- successors 1398 1402 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_trigger_
      -- 
    cpelement_group_1397 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1400);
      predecessors(1) <= cp_elements(1401);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1397)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1397),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1398 join  fork  transition  no-bypass 
    -- predecessors 1397 1403 
    -- successors 1399 1404 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_active_
      -- 
    cpelement_group_1398 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1397);
      predecessors(1) <= cp_elements(1403);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1398)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1398),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1399 join  transition  bypass 
    -- predecessors 1398 1405 
    -- successors 1406 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1327_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1327_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1327_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1330_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1330_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1330_completed_
      -- 
    cpelement_group_1399 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1398);
      predecessors(1) <= cp_elements(1405);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1399)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1399),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1400 transition  bypass 
    -- predecessors 1029 
    -- successors 1397 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1324_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1324_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1324_completed_
      -- 
    cp_elements(1400) <= cp_elements(1029);
    -- CP-element group 1401 transition  bypass 
    -- predecessors 1354 
    -- successors 1397 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1325_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1325_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1325_completed_
      -- 
    cp_elements(1401) <= cp_elements(1354);
    -- CP-element group 1402 transition  output  bypass 
    -- predecessors 1397 
    -- successors 1403 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Sample/rr
      -- 
    cp_elements(1402) <= cp_elements(1397);
    rr_6289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1402), ack => binary_1326_inst_req_0); -- 
    -- CP-element group 1403 transition  input  no-bypass 
    -- predecessors 1402 
    -- successors 1398 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Sample/ra
      -- 
    ra_6290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1326_inst_ack_0, ack => cp_elements(1403)); -- 
    -- CP-element group 1404 transition  output  bypass 
    -- predecessors 1398 
    -- successors 1405 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Update/cr
      -- 
    cp_elements(1404) <= cp_elements(1398);
    cr_6294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1404), ack => binary_1326_inst_req_1); -- 
    -- CP-element group 1405 transition  input  no-bypass 
    -- predecessors 1404 
    -- successors 1399 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1326_complete_Update/ca
      -- 
    ca_6295_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1326_inst_ack_1, ack => cp_elements(1405)); -- 
    -- CP-element group 1406 join  fork  transition  bypass 
    -- predecessors 1390 1399 
    -- successors 1407 1409 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_trigger_
      -- 
    cpelement_group_1406 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1390);
      predecessors(1) <= cp_elements(1399);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1406)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1406),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1407 join  fork  transition  no-bypass 
    -- predecessors 1406 1410 
    -- successors 1408 1411 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_active_
      -- 
    cpelement_group_1407 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1406);
      predecessors(1) <= cp_elements(1410);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1407)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1407),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1408 join  transition  no-bypass 
    -- predecessors 1407 1412 
    -- successors 1413 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1332_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1332_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1332_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1335_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1335_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1335_completed_
      -- 
    cpelement_group_1408 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1407);
      predecessors(1) <= cp_elements(1412);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1408)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1408),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1409 transition  output  bypass 
    -- predecessors 1406 
    -- successors 1410 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Sample/rr
      -- 
    cp_elements(1409) <= cp_elements(1406);
    rr_6311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1409), ack => binary_1331_inst_req_0); -- 
    -- CP-element group 1410 transition  input  no-bypass 
    -- predecessors 1409 
    -- successors 1407 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Sample/ra
      -- 
    ra_6312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1331_inst_ack_0, ack => cp_elements(1410)); -- 
    -- CP-element group 1411 transition  output  bypass 
    -- predecessors 1407 
    -- successors 1412 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Update/cr
      -- 
    cp_elements(1411) <= cp_elements(1407);
    cr_6316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1411), ack => binary_1331_inst_req_1); -- 
    -- CP-element group 1412 transition  input  no-bypass 
    -- predecessors 1411 
    -- successors 1408 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1331_complete_Update/ca
      -- 
    ca_6317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1331_inst_ack_1, ack => cp_elements(1412)); -- 
    -- CP-element group 1413 join  fork  transition  bypass 
    -- predecessors 1383 1408 
    -- successors 1414 1416 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_trigger_
      -- 
    cpelement_group_1413 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1383);
      predecessors(1) <= cp_elements(1408);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1413)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1413),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1414 join  fork  transition  no-bypass 
    -- predecessors 1413 1417 
    -- successors 1415 1418 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_active_
      -- 
    cpelement_group_1414 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1413);
      predecessors(1) <= cp_elements(1417);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1414)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1414),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1415 join  transition  no-bypass 
    -- predecessors 1414 1419 
    -- successors 1420 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1337_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1337_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1337_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1340_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1340_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1340_completed_
      -- 
    cpelement_group_1415 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1414);
      predecessors(1) <= cp_elements(1419);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1415)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1415),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1416 transition  output  bypass 
    -- predecessors 1413 
    -- successors 1417 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Sample/rr
      -- 
    cp_elements(1416) <= cp_elements(1413);
    rr_6333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1416), ack => binary_1336_inst_req_0); -- 
    -- CP-element group 1417 transition  input  no-bypass 
    -- predecessors 1416 
    -- successors 1414 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Sample/ra
      -- 
    ra_6334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1336_inst_ack_0, ack => cp_elements(1417)); -- 
    -- CP-element group 1418 transition  output  bypass 
    -- predecessors 1414 
    -- successors 1419 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Update/cr
      -- 
    cp_elements(1418) <= cp_elements(1414);
    cr_6338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1418), ack => binary_1336_inst_req_1); -- 
    -- CP-element group 1419 transition  input  no-bypass 
    -- predecessors 1418 
    -- successors 1415 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1336_complete_Update/ca
      -- 
    ca_6339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1336_inst_ack_1, ack => cp_elements(1419)); -- 
    -- CP-element group 1420 join  fork  transition  no-bypass 
    -- predecessors 1415 1423 
    -- successors 1421 1424 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_trigger_
      -- 
    cpelement_group_1420 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1415);
      predecessors(1) <= cp_elements(1423);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1420)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1420),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1421 join  fork  transition  bypass 
    -- predecessors 1420 1425 
    -- successors 1422 1426 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_active_
      -- 
    cpelement_group_1421 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1420);
      predecessors(1) <= cp_elements(1425);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1421)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1421),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1422 join  transition  bypass 
    -- predecessors 1421 1427 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1342_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1342_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1342_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_completed_
      -- 
    cpelement_group_1422 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1421);
      predecessors(1) <= cp_elements(1427);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1422)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1422),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1423 transition  bypass 
    -- predecessors 367 
    -- successors 1420 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1339_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1339_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1339_completed_
      -- 
    cp_elements(1423) <= cp_elements(367);
    -- CP-element group 1424 transition  output  bypass 
    -- predecessors 1420 
    -- successors 1425 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Sample/rr
      -- 
    cp_elements(1424) <= cp_elements(1420);
    rr_6355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1424), ack => binary_1341_inst_req_0); -- 
    -- CP-element group 1425 transition  input  no-bypass 
    -- predecessors 1424 
    -- successors 1421 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Sample/ra
      -- 
    ra_6356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1341_inst_ack_0, ack => cp_elements(1425)); -- 
    -- CP-element group 1426 transition  output  bypass 
    -- predecessors 1421 
    -- successors 1427 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Update/cr
      -- 
    cp_elements(1426) <= cp_elements(1421);
    cr_6360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1426), ack => binary_1341_inst_req_1); -- 
    -- CP-element group 1427 transition  input  no-bypass 
    -- predecessors 1426 
    -- successors 1422 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1341_complete_Update/ca
      -- 
    ca_6361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1341_inst_ack_1, ack => cp_elements(1427)); -- 
    -- CP-element group 1428 join  fork  transition  bypass 
    -- predecessors 1432 1434 
    -- successors 1429 1435 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_active_
      -- 
    cpelement_group_1428 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1432);
      predecessors(1) <= cp_elements(1434);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1428)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1428),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1429 join  fork  transition  bypass 
    -- predecessors 1428 1437 
    -- successors 1471 1536 1601 1666 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1346_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1346_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1346_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_completed_
      -- 
    cpelement_group_1429 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1428);
      predecessors(1) <= cp_elements(1437);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1429)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1429),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1430 transition  input  output  no-bypass 
    -- predecessors 585 
    -- successors 1431 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6379_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_base_resize_ack_0, ack => cp_elements(1430)); -- 
    sum_rename_req_6383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1430), ack => ptr_deref_1345_root_address_inst_req_0); -- 
    -- CP-element group 1431 transition  input  output  no-bypass 
    -- predecessors 1430 
    -- successors 1432 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_root_address_inst_ack_0, ack => cp_elements(1431)); -- 
    root_register_req_6388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1431), ack => ptr_deref_1345_addr_0_req_0); -- 
    -- CP-element group 1432 fork  transition  input  no-bypass 
    -- predecessors 1431 
    -- successors 1428 1433 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_word_addrgen/root_register_ack
      -- 
    root_register_ack_6389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_addr_0_ack_0, ack => cp_elements(1432)); -- 
    -- CP-element group 1433 transition  output  bypass 
    -- predecessors 1432 
    -- successors 1434 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/word_access/word_access_0/rr
      -- 
    cp_elements(1433) <= cp_elements(1432);
    rr_6399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1433), ack => ptr_deref_1345_load_0_req_0); -- 
    -- CP-element group 1434 transition  input  no-bypass 
    -- predecessors 1433 
    -- successors 1428 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_request/word_access/word_access_0/ra
      -- 
    ra_6400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_load_0_ack_0, ack => cp_elements(1434)); -- 
    -- CP-element group 1435 transition  output  bypass 
    -- predecessors 1428 
    -- successors 1436 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1435) <= cp_elements(1428);
    cr_6410_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1435), ack => ptr_deref_1345_load_0_req_1); -- 
    -- CP-element group 1436 transition  input  output  no-bypass 
    -- predecessors 1435 
    -- successors 1437 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/merge_req
      -- 
    ca_6411_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_load_0_ack_1, ack => cp_elements(1436)); -- 
    merge_req_6412_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1436), ack => ptr_deref_1345_gather_scatter_req_0); -- 
    -- CP-element group 1437 transition  input  no-bypass 
    -- predecessors 1436 
    -- successors 1429 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1345_complete/merge_ack
      -- 
    merge_ack_6413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_gather_scatter_ack_0, ack => cp_elements(1437)); -- 
    -- CP-element group 1438 join  fork  transition  bypass 
    -- predecessors 1442 1444 
    -- successors 1439 1445 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_active_
      -- 
    cpelement_group_1438 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1442);
      predecessors(1) <= cp_elements(1444);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1438)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1438),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1439 join  fork  transition  bypass 
    -- predecessors 1438 1447 
    -- successors 1480 1545 1610 1675 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1350_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1350_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1350_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_completed_
      -- 
    cpelement_group_1439 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1438);
      predecessors(1) <= cp_elements(1447);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1439)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1439),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1440 transition  input  output  no-bypass 
    -- predecessors 636 
    -- successors 1441 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1349_base_resize_ack_0, ack => cp_elements(1440)); -- 
    sum_rename_req_6435_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1440), ack => ptr_deref_1349_root_address_inst_req_0); -- 
    -- CP-element group 1441 transition  input  output  no-bypass 
    -- predecessors 1440 
    -- successors 1442 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6436_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1349_root_address_inst_ack_0, ack => cp_elements(1441)); -- 
    root_register_req_6440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1441), ack => ptr_deref_1349_addr_0_req_0); -- 
    -- CP-element group 1442 fork  transition  input  no-bypass 
    -- predecessors 1441 
    -- successors 1438 1443 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_word_addrgen/root_register_ack
      -- 
    root_register_ack_6441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1349_addr_0_ack_0, ack => cp_elements(1442)); -- 
    -- CP-element group 1443 transition  output  bypass 
    -- predecessors 1442 
    -- successors 1444 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/word_access/word_access_0/rr
      -- 
    cp_elements(1443) <= cp_elements(1442);
    rr_6451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1443), ack => ptr_deref_1349_load_0_req_0); -- 
    -- CP-element group 1444 transition  input  no-bypass 
    -- predecessors 1443 
    -- successors 1438 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_request/word_access/word_access_0/ra
      -- 
    ra_6452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1349_load_0_ack_0, ack => cp_elements(1444)); -- 
    -- CP-element group 1445 transition  output  bypass 
    -- predecessors 1438 
    -- successors 1446 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1445) <= cp_elements(1438);
    cr_6462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1445), ack => ptr_deref_1349_load_0_req_1); -- 
    -- CP-element group 1446 transition  input  output  no-bypass 
    -- predecessors 1445 
    -- successors 1447 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/merge_req
      -- 
    ca_6463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1349_load_0_ack_1, ack => cp_elements(1446)); -- 
    merge_req_6464_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1446), ack => ptr_deref_1349_gather_scatter_req_0); -- 
    -- CP-element group 1447 transition  input  no-bypass 
    -- predecessors 1446 
    -- successors 1439 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1349_complete/merge_ack
      -- 
    merge_ack_6465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1349_gather_scatter_ack_0, ack => cp_elements(1447)); -- 
    -- CP-element group 1448 join  fork  transition  bypass 
    -- predecessors 1452 1454 
    -- successors 1449 1455 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_active_
      -- 
    cpelement_group_1448 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1452);
      predecessors(1) <= cp_elements(1454);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1448)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1448),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1449 join  fork  transition  bypass 
    -- predecessors 1448 1457 
    -- successors 1496 1561 1626 1691 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1354_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1354_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1354_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_completed_
      -- 
    cpelement_group_1449 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1448);
      predecessors(1) <= cp_elements(1457);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1449)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1449),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1450 transition  input  output  no-bypass 
    -- predecessors 619 
    -- successors 1451 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_base_resize_ack_0, ack => cp_elements(1450)); -- 
    sum_rename_req_6487_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1450), ack => ptr_deref_1353_root_address_inst_req_0); -- 
    -- CP-element group 1451 transition  input  output  no-bypass 
    -- predecessors 1450 
    -- successors 1452 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6488_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_root_address_inst_ack_0, ack => cp_elements(1451)); -- 
    root_register_req_6492_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1451), ack => ptr_deref_1353_addr_0_req_0); -- 
    -- CP-element group 1452 fork  transition  input  no-bypass 
    -- predecessors 1451 
    -- successors 1448 1453 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_word_addrgen/root_register_ack
      -- 
    root_register_ack_6493_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_addr_0_ack_0, ack => cp_elements(1452)); -- 
    -- CP-element group 1453 transition  output  bypass 
    -- predecessors 1452 
    -- successors 1454 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/word_access/word_access_0/rr
      -- 
    cp_elements(1453) <= cp_elements(1452);
    rr_6503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1453), ack => ptr_deref_1353_load_0_req_0); -- 
    -- CP-element group 1454 transition  input  no-bypass 
    -- predecessors 1453 
    -- successors 1448 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_request/word_access/word_access_0/ra
      -- 
    ra_6504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_load_0_ack_0, ack => cp_elements(1454)); -- 
    -- CP-element group 1455 transition  output  bypass 
    -- predecessors 1448 
    -- successors 1456 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1455) <= cp_elements(1448);
    cr_6514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1455), ack => ptr_deref_1353_load_0_req_1); -- 
    -- CP-element group 1456 transition  input  output  no-bypass 
    -- predecessors 1455 
    -- successors 1457 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/merge_req
      -- 
    ca_6515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_load_0_ack_1, ack => cp_elements(1456)); -- 
    merge_req_6516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1456), ack => ptr_deref_1353_gather_scatter_req_0); -- 
    -- CP-element group 1457 transition  input  no-bypass 
    -- predecessors 1456 
    -- successors 1449 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1353_complete/merge_ack
      -- 
    merge_ack_6517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1353_gather_scatter_ack_0, ack => cp_elements(1457)); -- 
    -- CP-element group 1458 join  fork  transition  bypass 
    -- predecessors 1462 1464 
    -- successors 1459 1465 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_active_
      -- 
    cpelement_group_1458 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1462);
      predecessors(1) <= cp_elements(1464);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1458)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1458),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1459 join  fork  transition  bypass 
    -- predecessors 1458 1467 
    -- successors 1505 1570 1635 1700 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1358_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1358_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1358_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_completed_
      -- 
    cpelement_group_1459 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1458);
      predecessors(1) <= cp_elements(1467);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1459)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1459),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1460 transition  input  output  no-bypass 
    -- predecessors 602 
    -- successors 1461 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6535_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_base_resize_ack_0, ack => cp_elements(1460)); -- 
    sum_rename_req_6539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1460), ack => ptr_deref_1357_root_address_inst_req_0); -- 
    -- CP-element group 1461 transition  input  output  no-bypass 
    -- predecessors 1460 
    -- successors 1462 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_root_address_inst_ack_0, ack => cp_elements(1461)); -- 
    root_register_req_6544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1461), ack => ptr_deref_1357_addr_0_req_0); -- 
    -- CP-element group 1462 fork  transition  input  no-bypass 
    -- predecessors 1461 
    -- successors 1458 1463 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_word_addrgen/root_register_ack
      -- 
    root_register_ack_6545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_addr_0_ack_0, ack => cp_elements(1462)); -- 
    -- CP-element group 1463 transition  output  bypass 
    -- predecessors 1462 
    -- successors 1464 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/word_access/word_access_0/rr
      -- 
    cp_elements(1463) <= cp_elements(1462);
    rr_6555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1463), ack => ptr_deref_1357_load_0_req_0); -- 
    -- CP-element group 1464 transition  input  no-bypass 
    -- predecessors 1463 
    -- successors 1458 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_request/word_access/word_access_0/ra
      -- 
    ra_6556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_load_0_ack_0, ack => cp_elements(1464)); -- 
    -- CP-element group 1465 transition  output  bypass 
    -- predecessors 1458 
    -- successors 1466 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1465) <= cp_elements(1458);
    cr_6566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1465), ack => ptr_deref_1357_load_0_req_1); -- 
    -- CP-element group 1466 transition  input  output  no-bypass 
    -- predecessors 1465 
    -- successors 1467 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/merge_req
      -- 
    ca_6567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_load_0_ack_1, ack => cp_elements(1466)); -- 
    merge_req_6568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1466), ack => ptr_deref_1357_gather_scatter_req_0); -- 
    -- CP-element group 1467 transition  input  no-bypass 
    -- predecessors 1466 
    -- successors 1459 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1357_complete/merge_ack
      -- 
    merge_ack_6569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_gather_scatter_ack_0, ack => cp_elements(1467)); -- 
    -- CP-element group 1468 join  fork  transition  no-bypass 
    -- predecessors 1471 1472 
    -- successors 1469 1473 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_trigger_
      -- 
    cpelement_group_1468 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1471);
      predecessors(1) <= cp_elements(1472);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1468)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1468),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1469 join  fork  transition  no-bypass 
    -- predecessors 1468 1474 
    -- successors 1470 1475 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_active_
      -- 
    cpelement_group_1469 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1468);
      predecessors(1) <= cp_elements(1474);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1469)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1469),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1470 join  transition  bypass 
    -- predecessors 1469 1476 
    -- successors 1486 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1363_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1363_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1363_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1370_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1370_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1370_completed_
      -- 
    cpelement_group_1470 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1469);
      predecessors(1) <= cp_elements(1476);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1470)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1470),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1471 transition  bypass 
    -- predecessors 1429 
    -- successors 1468 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1360_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1360_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1360_completed_
      -- 
    cp_elements(1471) <= cp_elements(1429);
    -- CP-element group 1472 transition  bypass 
    -- predecessors 979 
    -- successors 1468 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1361_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1361_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1361_completed_
      -- 
    cp_elements(1472) <= cp_elements(979);
    -- CP-element group 1473 transition  output  bypass 
    -- predecessors 1468 
    -- successors 1474 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Sample/rr
      -- 
    cp_elements(1473) <= cp_elements(1468);
    rr_6585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1473), ack => binary_1362_inst_req_0); -- 
    -- CP-element group 1474 transition  input  no-bypass 
    -- predecessors 1473 
    -- successors 1469 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Sample/ra
      -- 
    ra_6586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1362_inst_ack_0, ack => cp_elements(1474)); -- 
    -- CP-element group 1475 transition  output  bypass 
    -- predecessors 1469 
    -- successors 1476 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Update/cr
      -- 
    cp_elements(1475) <= cp_elements(1469);
    cr_6590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1475), ack => binary_1362_inst_req_1); -- 
    -- CP-element group 1476 transition  input  no-bypass 
    -- predecessors 1475 
    -- successors 1470 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1362_complete_Update/ca
      -- 
    ca_6591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1362_inst_ack_1, ack => cp_elements(1476)); -- 
    -- CP-element group 1477 join  fork  transition  no-bypass 
    -- predecessors 1480 1481 
    -- successors 1478 1482 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_trigger_
      -- 
    cpelement_group_1477 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1480);
      predecessors(1) <= cp_elements(1481);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1477)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1477),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1478 join  fork  transition  no-bypass 
    -- predecessors 1477 1483 
    -- successors 1479 1484 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_active_
      -- 
    cpelement_group_1478 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1477);
      predecessors(1) <= cp_elements(1483);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1478)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1478),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1479 join  transition  bypass 
    -- predecessors 1478 1485 
    -- successors 1486 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1368_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1368_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1368_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1371_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1371_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1371_completed_
      -- 
    cpelement_group_1479 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1478);
      predecessors(1) <= cp_elements(1485);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1479)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1479),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1480 transition  bypass 
    -- predecessors 1439 
    -- successors 1477 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1365_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1365_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1365_completed_
      -- 
    cp_elements(1480) <= cp_elements(1439);
    -- CP-element group 1481 transition  bypass 
    -- predecessors 999 
    -- successors 1477 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1366_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1366_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1366_completed_
      -- 
    cp_elements(1481) <= cp_elements(999);
    -- CP-element group 1482 transition  output  bypass 
    -- predecessors 1477 
    -- successors 1483 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Sample/rr
      -- 
    cp_elements(1482) <= cp_elements(1477);
    rr_6607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1482), ack => binary_1367_inst_req_0); -- 
    -- CP-element group 1483 transition  input  no-bypass 
    -- predecessors 1482 
    -- successors 1478 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Sample/ra
      -- 
    ra_6608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1367_inst_ack_0, ack => cp_elements(1483)); -- 
    -- CP-element group 1484 transition  output  bypass 
    -- predecessors 1478 
    -- successors 1485 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Update/cr
      -- 
    cp_elements(1484) <= cp_elements(1478);
    cr_6612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1484), ack => binary_1367_inst_req_1); -- 
    -- CP-element group 1485 transition  input  no-bypass 
    -- predecessors 1484 
    -- successors 1479 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1367_complete_Update/ca
      -- 
    ca_6613_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1367_inst_ack_1, ack => cp_elements(1485)); -- 
    -- CP-element group 1486 join  fork  transition  bypass 
    -- predecessors 1470 1479 
    -- successors 1487 1489 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_trigger_
      -- 
    cpelement_group_1486 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1470);
      predecessors(1) <= cp_elements(1479);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1486)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1486),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1487 join  fork  transition  no-bypass 
    -- predecessors 1486 1490 
    -- successors 1488 1491 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_active_
      -- 
    cpelement_group_1487 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1486);
      predecessors(1) <= cp_elements(1490);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1487)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1487),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1488 join  transition  no-bypass 
    -- predecessors 1487 1492 
    -- successors 1518 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1373_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1373_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1373_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1390_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1390_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1390_completed_
      -- 
    cpelement_group_1488 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1487);
      predecessors(1) <= cp_elements(1492);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1488)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1488),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1489 transition  output  bypass 
    -- predecessors 1486 
    -- successors 1490 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Sample/rr
      -- 
    cp_elements(1489) <= cp_elements(1486);
    rr_6629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1489), ack => binary_1372_inst_req_0); -- 
    -- CP-element group 1490 transition  input  no-bypass 
    -- predecessors 1489 
    -- successors 1487 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Sample/ra
      -- 
    ra_6630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1372_inst_ack_0, ack => cp_elements(1490)); -- 
    -- CP-element group 1491 transition  output  bypass 
    -- predecessors 1487 
    -- successors 1492 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Update/cr
      -- 
    cp_elements(1491) <= cp_elements(1487);
    cr_6634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1491), ack => binary_1372_inst_req_1); -- 
    -- CP-element group 1492 transition  input  no-bypass 
    -- predecessors 1491 
    -- successors 1488 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1372_complete_Update/ca
      -- 
    ca_6635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1372_inst_ack_1, ack => cp_elements(1492)); -- 
    -- CP-element group 1493 join  fork  transition  no-bypass 
    -- predecessors 1496 1497 
    -- successors 1494 1498 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_trigger_
      -- 
    cpelement_group_1493 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1496);
      predecessors(1) <= cp_elements(1497);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1493)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1493),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1494 join  fork  transition  no-bypass 
    -- predecessors 1493 1499 
    -- successors 1495 1500 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_active_
      -- 
    cpelement_group_1494 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1493);
      predecessors(1) <= cp_elements(1499);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1494)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1494),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1495 join  transition  bypass 
    -- predecessors 1494 1501 
    -- successors 1511 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1378_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1378_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1378_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1385_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1385_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1385_completed_
      -- 
    cpelement_group_1495 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1494);
      predecessors(1) <= cp_elements(1501);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1495)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1495),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1496 transition  bypass 
    -- predecessors 1449 
    -- successors 1493 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1375_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1375_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1375_completed_
      -- 
    cp_elements(1496) <= cp_elements(1449);
    -- CP-element group 1497 transition  bypass 
    -- predecessors 1019 
    -- successors 1493 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1376_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1376_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1376_completed_
      -- 
    cp_elements(1497) <= cp_elements(1019);
    -- CP-element group 1498 transition  output  bypass 
    -- predecessors 1493 
    -- successors 1499 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Sample/rr
      -- 
    cp_elements(1498) <= cp_elements(1493);
    rr_6651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1498), ack => binary_1377_inst_req_0); -- 
    -- CP-element group 1499 transition  input  no-bypass 
    -- predecessors 1498 
    -- successors 1494 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Sample/ra
      -- 
    ra_6652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1377_inst_ack_0, ack => cp_elements(1499)); -- 
    -- CP-element group 1500 transition  output  bypass 
    -- predecessors 1494 
    -- successors 1501 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Update/cr
      -- 
    cp_elements(1500) <= cp_elements(1494);
    cr_6656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1500), ack => binary_1377_inst_req_1); -- 
    -- CP-element group 1501 transition  input  no-bypass 
    -- predecessors 1500 
    -- successors 1495 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1377_complete_Update/ca
      -- 
    ca_6657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1377_inst_ack_1, ack => cp_elements(1501)); -- 
    -- CP-element group 1502 join  fork  transition  no-bypass 
    -- predecessors 1505 1506 
    -- successors 1503 1507 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_trigger_
      -- 
    cpelement_group_1502 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1505);
      predecessors(1) <= cp_elements(1506);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1502)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1502),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1503 join  fork  transition  no-bypass 
    -- predecessors 1502 1508 
    -- successors 1504 1509 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_active_
      -- 
    cpelement_group_1503 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1502);
      predecessors(1) <= cp_elements(1508);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1503)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1503),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1504 join  transition  bypass 
    -- predecessors 1503 1510 
    -- successors 1511 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1383_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1383_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1383_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1386_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1386_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1386_completed_
      -- 
    cpelement_group_1504 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1503);
      predecessors(1) <= cp_elements(1510);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1504)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1504),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1505 transition  bypass 
    -- predecessors 1459 
    -- successors 1502 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1380_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1380_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1380_completed_
      -- 
    cp_elements(1505) <= cp_elements(1459);
    -- CP-element group 1506 transition  bypass 
    -- predecessors 1039 
    -- successors 1502 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1381_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1381_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1381_completed_
      -- 
    cp_elements(1506) <= cp_elements(1039);
    -- CP-element group 1507 transition  output  bypass 
    -- predecessors 1502 
    -- successors 1508 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Sample/rr
      -- 
    cp_elements(1507) <= cp_elements(1502);
    rr_6673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1507), ack => binary_1382_inst_req_0); -- 
    -- CP-element group 1508 transition  input  no-bypass 
    -- predecessors 1507 
    -- successors 1503 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Sample/ra
      -- 
    ra_6674_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1382_inst_ack_0, ack => cp_elements(1508)); -- 
    -- CP-element group 1509 transition  output  bypass 
    -- predecessors 1503 
    -- successors 1510 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Update/cr
      -- 
    cp_elements(1509) <= cp_elements(1503);
    cr_6678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1509), ack => binary_1382_inst_req_1); -- 
    -- CP-element group 1510 transition  input  no-bypass 
    -- predecessors 1509 
    -- successors 1504 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1382_complete_Update/ca
      -- 
    ca_6679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1382_inst_ack_1, ack => cp_elements(1510)); -- 
    -- CP-element group 1511 join  fork  transition  bypass 
    -- predecessors 1495 1504 
    -- successors 1512 1514 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_trigger_
      -- 
    cpelement_group_1511 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1495);
      predecessors(1) <= cp_elements(1504);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1511)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1511),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1512 join  fork  transition  no-bypass 
    -- predecessors 1511 1515 
    -- successors 1513 1516 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_active_
      -- 
    cpelement_group_1512 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1511);
      predecessors(1) <= cp_elements(1515);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1512)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1512),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1513 join  transition  no-bypass 
    -- predecessors 1512 1517 
    -- successors 1518 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1388_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1388_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1388_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1391_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1391_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1391_completed_
      -- 
    cpelement_group_1513 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1512);
      predecessors(1) <= cp_elements(1517);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1513)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1513),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1514 transition  output  bypass 
    -- predecessors 1511 
    -- successors 1515 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Sample/rr
      -- 
    cp_elements(1514) <= cp_elements(1511);
    rr_6695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1514), ack => binary_1387_inst_req_0); -- 
    -- CP-element group 1515 transition  input  no-bypass 
    -- predecessors 1514 
    -- successors 1512 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Sample/ra
      -- 
    ra_6696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1387_inst_ack_0, ack => cp_elements(1515)); -- 
    -- CP-element group 1516 transition  output  bypass 
    -- predecessors 1512 
    -- successors 1517 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Update/cr
      -- 
    cp_elements(1516) <= cp_elements(1512);
    cr_6700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1516), ack => binary_1387_inst_req_1); -- 
    -- CP-element group 1517 transition  input  no-bypass 
    -- predecessors 1516 
    -- successors 1513 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1387_complete_Update/ca
      -- 
    ca_6701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1387_inst_ack_1, ack => cp_elements(1517)); -- 
    -- CP-element group 1518 join  fork  transition  bypass 
    -- predecessors 1488 1513 
    -- successors 1519 1521 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_trigger_
      -- 
    cpelement_group_1518 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1488);
      predecessors(1) <= cp_elements(1513);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1518)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1518),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1519 join  fork  transition  no-bypass 
    -- predecessors 1518 1522 
    -- successors 1520 1523 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_active_
      -- 
    cpelement_group_1519 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1518);
      predecessors(1) <= cp_elements(1522);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1519)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1519),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1520 join  transition  no-bypass 
    -- predecessors 1519 1524 
    -- successors 1525 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1393_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1393_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1393_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1396_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1396_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1396_completed_
      -- 
    cpelement_group_1520 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1519);
      predecessors(1) <= cp_elements(1524);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1520)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1520),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1521 transition  output  bypass 
    -- predecessors 1518 
    -- successors 1522 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Sample/rr
      -- 
    cp_elements(1521) <= cp_elements(1518);
    rr_6717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1521), ack => binary_1392_inst_req_0); -- 
    -- CP-element group 1522 transition  input  no-bypass 
    -- predecessors 1521 
    -- successors 1519 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Sample/ra
      -- 
    ra_6718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1392_inst_ack_0, ack => cp_elements(1522)); -- 
    -- CP-element group 1523 transition  output  bypass 
    -- predecessors 1519 
    -- successors 1524 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Update/cr
      -- 
    cp_elements(1523) <= cp_elements(1519);
    cr_6722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1523), ack => binary_1392_inst_req_1); -- 
    -- CP-element group 1524 transition  input  no-bypass 
    -- predecessors 1523 
    -- successors 1520 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1392_complete_Update/ca
      -- 
    ca_6723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1392_inst_ack_1, ack => cp_elements(1524)); -- 
    -- CP-element group 1525 join  fork  transition  no-bypass 
    -- predecessors 1520 1528 
    -- successors 1526 1529 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_trigger_
      -- 
    cpelement_group_1525 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1520);
      predecessors(1) <= cp_elements(1528);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1525)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1525),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1526 join  fork  transition  bypass 
    -- predecessors 1525 1530 
    -- successors 1527 1531 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_active_
      -- 
    cpelement_group_1526 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1525);
      predecessors(1) <= cp_elements(1530);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1526)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1526),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1527 join  transition  bypass 
    -- predecessors 1526 1532 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1398_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1398_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1398_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_completed_
      -- 
    cpelement_group_1527 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1526);
      predecessors(1) <= cp_elements(1532);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1527)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1527),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1528 transition  bypass 
    -- predecessors 367 
    -- successors 1525 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1395_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1395_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1395_completed_
      -- 
    cp_elements(1528) <= cp_elements(367);
    -- CP-element group 1529 transition  output  bypass 
    -- predecessors 1525 
    -- successors 1530 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Sample/rr
      -- 
    cp_elements(1529) <= cp_elements(1525);
    rr_6739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1529), ack => binary_1397_inst_req_0); -- 
    -- CP-element group 1530 transition  input  no-bypass 
    -- predecessors 1529 
    -- successors 1526 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Sample/ra
      -- 
    ra_6740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1397_inst_ack_0, ack => cp_elements(1530)); -- 
    -- CP-element group 1531 transition  output  bypass 
    -- predecessors 1526 
    -- successors 1532 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Update/cr
      -- 
    cp_elements(1531) <= cp_elements(1526);
    cr_6744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1531), ack => binary_1397_inst_req_1); -- 
    -- CP-element group 1532 transition  input  no-bypass 
    -- predecessors 1531 
    -- successors 1527 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1397_complete_Update/ca
      -- 
    ca_6745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1397_inst_ack_1, ack => cp_elements(1532)); -- 
    -- CP-element group 1533 join  fork  transition  no-bypass 
    -- predecessors 1536 1537 
    -- successors 1534 1538 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_trigger_
      -- 
    cpelement_group_1533 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1536);
      predecessors(1) <= cp_elements(1537);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1533)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1533),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1534 join  fork  transition  no-bypass 
    -- predecessors 1533 1539 
    -- successors 1535 1540 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_active_
      -- 
    cpelement_group_1534 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1533);
      predecessors(1) <= cp_elements(1539);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1534)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1534),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1535 join  transition  bypass 
    -- predecessors 1534 1541 
    -- successors 1551 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1403_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1403_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1403_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1410_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1410_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1410_completed_
      -- 
    cpelement_group_1535 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1534);
      predecessors(1) <= cp_elements(1541);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1535)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1535),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1536 transition  bypass 
    -- predecessors 1429 
    -- successors 1533 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1400_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1400_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1400_completed_
      -- 
    cp_elements(1536) <= cp_elements(1429);
    -- CP-element group 1537 transition  bypass 
    -- predecessors 1114 
    -- successors 1533 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1401_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1401_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1401_completed_
      -- 
    cp_elements(1537) <= cp_elements(1114);
    -- CP-element group 1538 transition  output  bypass 
    -- predecessors 1533 
    -- successors 1539 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Sample/rr
      -- 
    cp_elements(1538) <= cp_elements(1533);
    rr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1538), ack => binary_1402_inst_req_0); -- 
    -- CP-element group 1539 transition  input  no-bypass 
    -- predecessors 1538 
    -- successors 1534 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Sample/ra
      -- 
    ra_6762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1402_inst_ack_0, ack => cp_elements(1539)); -- 
    -- CP-element group 1540 transition  output  bypass 
    -- predecessors 1534 
    -- successors 1541 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Update/cr
      -- 
    cp_elements(1540) <= cp_elements(1534);
    cr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1540), ack => binary_1402_inst_req_1); -- 
    -- CP-element group 1541 transition  input  no-bypass 
    -- predecessors 1540 
    -- successors 1535 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1402_complete_Update/ca
      -- 
    ca_6767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1402_inst_ack_1, ack => cp_elements(1541)); -- 
    -- CP-element group 1542 join  fork  transition  no-bypass 
    -- predecessors 1545 1546 
    -- successors 1543 1547 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_trigger_
      -- 
    cpelement_group_1542 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1545);
      predecessors(1) <= cp_elements(1546);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1542)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1542),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1543 join  fork  transition  no-bypass 
    -- predecessors 1542 1548 
    -- successors 1544 1549 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_active_
      -- 
    cpelement_group_1543 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1542);
      predecessors(1) <= cp_elements(1548);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1543)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1543),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1544 join  transition  bypass 
    -- predecessors 1543 1550 
    -- successors 1551 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1408_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1408_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1408_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1411_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1411_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1411_completed_
      -- 
    cpelement_group_1544 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1543);
      predecessors(1) <= cp_elements(1550);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1544)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1544),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1545 transition  bypass 
    -- predecessors 1439 
    -- successors 1542 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1405_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1405_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1405_completed_
      -- 
    cp_elements(1545) <= cp_elements(1439);
    -- CP-element group 1546 transition  bypass 
    -- predecessors 1124 
    -- successors 1542 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1406_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1406_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1406_completed_
      -- 
    cp_elements(1546) <= cp_elements(1124);
    -- CP-element group 1547 transition  output  bypass 
    -- predecessors 1542 
    -- successors 1548 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Sample/rr
      -- 
    cp_elements(1547) <= cp_elements(1542);
    rr_6783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1547), ack => binary_1407_inst_req_0); -- 
    -- CP-element group 1548 transition  input  no-bypass 
    -- predecessors 1547 
    -- successors 1543 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Sample/ra
      -- 
    ra_6784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1407_inst_ack_0, ack => cp_elements(1548)); -- 
    -- CP-element group 1549 transition  output  bypass 
    -- predecessors 1543 
    -- successors 1550 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Update/cr
      -- 
    cp_elements(1549) <= cp_elements(1543);
    cr_6788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1549), ack => binary_1407_inst_req_1); -- 
    -- CP-element group 1550 transition  input  no-bypass 
    -- predecessors 1549 
    -- successors 1544 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1407_complete_Update/ca
      -- 
    ca_6789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1407_inst_ack_1, ack => cp_elements(1550)); -- 
    -- CP-element group 1551 join  fork  transition  bypass 
    -- predecessors 1535 1544 
    -- successors 1552 1554 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_trigger_
      -- 
    cpelement_group_1551 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1535);
      predecessors(1) <= cp_elements(1544);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1551)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1551),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1552 join  fork  transition  no-bypass 
    -- predecessors 1551 1555 
    -- successors 1553 1556 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_active_
      -- 
    cpelement_group_1552 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1551);
      predecessors(1) <= cp_elements(1555);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1552)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1552),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1553 join  transition  no-bypass 
    -- predecessors 1552 1557 
    -- successors 1583 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1413_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1413_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1413_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1430_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1430_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1430_completed_
      -- 
    cpelement_group_1553 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1552);
      predecessors(1) <= cp_elements(1557);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1553)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1553),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1554 transition  output  bypass 
    -- predecessors 1551 
    -- successors 1555 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Sample/rr
      -- 
    cp_elements(1554) <= cp_elements(1551);
    rr_6805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1554), ack => binary_1412_inst_req_0); -- 
    -- CP-element group 1555 transition  input  no-bypass 
    -- predecessors 1554 
    -- successors 1552 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Sample/ra
      -- 
    ra_6806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1412_inst_ack_0, ack => cp_elements(1555)); -- 
    -- CP-element group 1556 transition  output  bypass 
    -- predecessors 1552 
    -- successors 1557 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Update/cr
      -- 
    cp_elements(1556) <= cp_elements(1552);
    cr_6810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1556), ack => binary_1412_inst_req_1); -- 
    -- CP-element group 1557 transition  input  no-bypass 
    -- predecessors 1556 
    -- successors 1553 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1412_complete_Update/ca
      -- 
    ca_6811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1412_inst_ack_1, ack => cp_elements(1557)); -- 
    -- CP-element group 1558 join  fork  transition  no-bypass 
    -- predecessors 1561 1562 
    -- successors 1559 1563 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_trigger_
      -- 
    cpelement_group_1558 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1561);
      predecessors(1) <= cp_elements(1562);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1558)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1558),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1559 join  fork  transition  no-bypass 
    -- predecessors 1558 1564 
    -- successors 1560 1565 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_active_
      -- 
    cpelement_group_1559 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1558);
      predecessors(1) <= cp_elements(1564);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1559)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1559),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1560 join  transition  bypass 
    -- predecessors 1559 1566 
    -- successors 1576 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1418_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1418_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1418_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1425_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1425_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1425_completed_
      -- 
    cpelement_group_1560 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1559);
      predecessors(1) <= cp_elements(1566);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1560)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1560),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1561 transition  bypass 
    -- predecessors 1449 
    -- successors 1558 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1415_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1415_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1415_completed_
      -- 
    cp_elements(1561) <= cp_elements(1449);
    -- CP-element group 1562 transition  bypass 
    -- predecessors 1134 
    -- successors 1558 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1416_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1416_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1416_completed_
      -- 
    cp_elements(1562) <= cp_elements(1134);
    -- CP-element group 1563 transition  output  bypass 
    -- predecessors 1558 
    -- successors 1564 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Sample/rr
      -- 
    cp_elements(1563) <= cp_elements(1558);
    rr_6827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1563), ack => binary_1417_inst_req_0); -- 
    -- CP-element group 1564 transition  input  no-bypass 
    -- predecessors 1563 
    -- successors 1559 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Sample/ra
      -- 
    ra_6828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1417_inst_ack_0, ack => cp_elements(1564)); -- 
    -- CP-element group 1565 transition  output  bypass 
    -- predecessors 1559 
    -- successors 1566 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Update/cr
      -- 
    cp_elements(1565) <= cp_elements(1559);
    cr_6832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1565), ack => binary_1417_inst_req_1); -- 
    -- CP-element group 1566 transition  input  no-bypass 
    -- predecessors 1565 
    -- successors 1560 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1417_complete_Update/ca
      -- 
    ca_6833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1417_inst_ack_1, ack => cp_elements(1566)); -- 
    -- CP-element group 1567 join  fork  transition  no-bypass 
    -- predecessors 1570 1571 
    -- successors 1568 1572 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_trigger_
      -- 
    cpelement_group_1567 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1570);
      predecessors(1) <= cp_elements(1571);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1567)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1567),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1568 join  fork  transition  no-bypass 
    -- predecessors 1567 1573 
    -- successors 1569 1574 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_active_
      -- 
    cpelement_group_1568 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1567);
      predecessors(1) <= cp_elements(1573);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1568)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1568),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1569 join  transition  bypass 
    -- predecessors 1568 1575 
    -- successors 1576 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1423_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1423_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1423_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1426_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1426_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1426_completed_
      -- 
    cpelement_group_1569 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1568);
      predecessors(1) <= cp_elements(1575);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1569)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1569),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1570 transition  bypass 
    -- predecessors 1459 
    -- successors 1567 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1420_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1420_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1420_completed_
      -- 
    cp_elements(1570) <= cp_elements(1459);
    -- CP-element group 1571 transition  bypass 
    -- predecessors 1144 
    -- successors 1567 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1421_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1421_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1421_completed_
      -- 
    cp_elements(1571) <= cp_elements(1144);
    -- CP-element group 1572 transition  output  bypass 
    -- predecessors 1567 
    -- successors 1573 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Sample/rr
      -- 
    cp_elements(1572) <= cp_elements(1567);
    rr_6849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1572), ack => binary_1422_inst_req_0); -- 
    -- CP-element group 1573 transition  input  no-bypass 
    -- predecessors 1572 
    -- successors 1568 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Sample/ra
      -- 
    ra_6850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1422_inst_ack_0, ack => cp_elements(1573)); -- 
    -- CP-element group 1574 transition  output  bypass 
    -- predecessors 1568 
    -- successors 1575 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Update/cr
      -- 
    cp_elements(1574) <= cp_elements(1568);
    cr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1574), ack => binary_1422_inst_req_1); -- 
    -- CP-element group 1575 transition  input  no-bypass 
    -- predecessors 1574 
    -- successors 1569 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1422_complete_Update/ca
      -- 
    ca_6855_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1422_inst_ack_1, ack => cp_elements(1575)); -- 
    -- CP-element group 1576 join  fork  transition  bypass 
    -- predecessors 1560 1569 
    -- successors 1577 1579 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_trigger_
      -- 
    cpelement_group_1576 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1560);
      predecessors(1) <= cp_elements(1569);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1576)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1576),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1577 join  fork  transition  no-bypass 
    -- predecessors 1576 1580 
    -- successors 1578 1581 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_active_
      -- 
    cpelement_group_1577 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1576);
      predecessors(1) <= cp_elements(1580);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1577)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1577),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1578 join  transition  no-bypass 
    -- predecessors 1577 1582 
    -- successors 1583 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1428_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1428_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1428_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1431_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1431_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1431_completed_
      -- 
    cpelement_group_1578 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1577);
      predecessors(1) <= cp_elements(1582);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1578)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1578),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1579 transition  output  bypass 
    -- predecessors 1576 
    -- successors 1580 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Sample/rr
      -- 
    cp_elements(1579) <= cp_elements(1576);
    rr_6871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1579), ack => binary_1427_inst_req_0); -- 
    -- CP-element group 1580 transition  input  no-bypass 
    -- predecessors 1579 
    -- successors 1577 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Sample/ra
      -- 
    ra_6872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1427_inst_ack_0, ack => cp_elements(1580)); -- 
    -- CP-element group 1581 transition  output  bypass 
    -- predecessors 1577 
    -- successors 1582 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Update/cr
      -- 
    cp_elements(1581) <= cp_elements(1577);
    cr_6876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1581), ack => binary_1427_inst_req_1); -- 
    -- CP-element group 1582 transition  input  no-bypass 
    -- predecessors 1581 
    -- successors 1578 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1427_complete_Update/ca
      -- 
    ca_6877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1427_inst_ack_1, ack => cp_elements(1582)); -- 
    -- CP-element group 1583 join  fork  transition  bypass 
    -- predecessors 1553 1578 
    -- successors 1584 1586 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_trigger_
      -- 
    cpelement_group_1583 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1553);
      predecessors(1) <= cp_elements(1578);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1583)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1583),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1584 join  fork  transition  no-bypass 
    -- predecessors 1583 1587 
    -- successors 1585 1588 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_active_
      -- 
    cpelement_group_1584 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1583);
      predecessors(1) <= cp_elements(1587);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1584)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1584),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1585 join  transition  no-bypass 
    -- predecessors 1584 1589 
    -- successors 1590 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1433_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1433_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1433_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1436_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1436_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1436_completed_
      -- 
    cpelement_group_1585 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1584);
      predecessors(1) <= cp_elements(1589);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1585)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1585),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1586 transition  output  bypass 
    -- predecessors 1583 
    -- successors 1587 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Sample/rr
      -- 
    cp_elements(1586) <= cp_elements(1583);
    rr_6893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1586), ack => binary_1432_inst_req_0); -- 
    -- CP-element group 1587 transition  input  no-bypass 
    -- predecessors 1586 
    -- successors 1584 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Sample/ra
      -- 
    ra_6894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1432_inst_ack_0, ack => cp_elements(1587)); -- 
    -- CP-element group 1588 transition  output  bypass 
    -- predecessors 1584 
    -- successors 1589 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Update/cr
      -- 
    cp_elements(1588) <= cp_elements(1584);
    cr_6898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1588), ack => binary_1432_inst_req_1); -- 
    -- CP-element group 1589 transition  input  no-bypass 
    -- predecessors 1588 
    -- successors 1585 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1432_complete_Update/ca
      -- 
    ca_6899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1432_inst_ack_1, ack => cp_elements(1589)); -- 
    -- CP-element group 1590 join  fork  transition  no-bypass 
    -- predecessors 1585 1593 
    -- successors 1591 1594 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_trigger_
      -- 
    cpelement_group_1590 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1585);
      predecessors(1) <= cp_elements(1593);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1590)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1590),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1591 join  fork  transition  bypass 
    -- predecessors 1590 1595 
    -- successors 1592 1596 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_active_
      -- 
    cpelement_group_1591 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1590);
      predecessors(1) <= cp_elements(1595);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1591)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1591),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1592 join  transition  bypass 
    -- predecessors 1591 1597 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1438_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1438_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1438_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_completed_
      -- 
    cpelement_group_1592 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1591);
      predecessors(1) <= cp_elements(1597);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1592)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1592),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1593 transition  bypass 
    -- predecessors 367 
    -- successors 1590 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1435_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1435_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1435_completed_
      -- 
    cp_elements(1593) <= cp_elements(367);
    -- CP-element group 1594 transition  output  bypass 
    -- predecessors 1590 
    -- successors 1595 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Sample/rr
      -- 
    cp_elements(1594) <= cp_elements(1590);
    rr_6915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1594), ack => binary_1437_inst_req_0); -- 
    -- CP-element group 1595 transition  input  no-bypass 
    -- predecessors 1594 
    -- successors 1591 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Sample/ra
      -- 
    ra_6916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1437_inst_ack_0, ack => cp_elements(1595)); -- 
    -- CP-element group 1596 transition  output  bypass 
    -- predecessors 1591 
    -- successors 1597 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Update/cr
      -- 
    cp_elements(1596) <= cp_elements(1591);
    cr_6920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1596), ack => binary_1437_inst_req_1); -- 
    -- CP-element group 1597 transition  input  no-bypass 
    -- predecessors 1596 
    -- successors 1592 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1437_complete_Update/ca
      -- 
    ca_6921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1437_inst_ack_1, ack => cp_elements(1597)); -- 
    -- CP-element group 1598 join  fork  transition  no-bypass 
    -- predecessors 1601 1602 
    -- successors 1599 1603 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_trigger_
      -- 
    cpelement_group_1598 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1601);
      predecessors(1) <= cp_elements(1602);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1598)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1598),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1599 join  fork  transition  no-bypass 
    -- predecessors 1598 1604 
    -- successors 1600 1605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_active_
      -- 
    cpelement_group_1599 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1598);
      predecessors(1) <= cp_elements(1604);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1599)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1599),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1600 join  transition  bypass 
    -- predecessors 1599 1606 
    -- successors 1616 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1443_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1443_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1443_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1450_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1450_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1450_completed_
      -- 
    cpelement_group_1600 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1599);
      predecessors(1) <= cp_elements(1606);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1600)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1600),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1601 transition  bypass 
    -- predecessors 1429 
    -- successors 1598 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1440_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1440_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1440_completed_
      -- 
    cp_elements(1601) <= cp_elements(1429);
    -- CP-element group 1602 transition  bypass 
    -- predecessors 1219 
    -- successors 1598 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1441_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1441_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1441_completed_
      -- 
    cp_elements(1602) <= cp_elements(1219);
    -- CP-element group 1603 transition  output  bypass 
    -- predecessors 1598 
    -- successors 1604 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Sample/rr
      -- 
    cp_elements(1603) <= cp_elements(1598);
    rr_6937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1603), ack => binary_1442_inst_req_0); -- 
    -- CP-element group 1604 transition  input  no-bypass 
    -- predecessors 1603 
    -- successors 1599 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Sample/ra
      -- 
    ra_6938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1442_inst_ack_0, ack => cp_elements(1604)); -- 
    -- CP-element group 1605 transition  output  bypass 
    -- predecessors 1599 
    -- successors 1606 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Update/cr
      -- 
    cp_elements(1605) <= cp_elements(1599);
    cr_6942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1605), ack => binary_1442_inst_req_1); -- 
    -- CP-element group 1606 transition  input  no-bypass 
    -- predecessors 1605 
    -- successors 1600 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1442_complete_Update/ca
      -- 
    ca_6943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1442_inst_ack_1, ack => cp_elements(1606)); -- 
    -- CP-element group 1607 join  fork  transition  no-bypass 
    -- predecessors 1610 1611 
    -- successors 1608 1612 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_trigger_
      -- 
    cpelement_group_1607 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1610);
      predecessors(1) <= cp_elements(1611);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1607)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1607),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1608 join  fork  transition  no-bypass 
    -- predecessors 1607 1613 
    -- successors 1609 1614 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_active_
      -- 
    cpelement_group_1608 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1607);
      predecessors(1) <= cp_elements(1613);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1608)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1608),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1609 join  transition  bypass 
    -- predecessors 1608 1615 
    -- successors 1616 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1448_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1448_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1448_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1451_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1451_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1451_completed_
      -- 
    cpelement_group_1609 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1608);
      predecessors(1) <= cp_elements(1615);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1609)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1609),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1610 transition  bypass 
    -- predecessors 1439 
    -- successors 1607 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1445_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1445_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1445_completed_
      -- 
    cp_elements(1610) <= cp_elements(1439);
    -- CP-element group 1611 transition  bypass 
    -- predecessors 1229 
    -- successors 1607 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1446_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1446_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1446_active_
      -- 
    cp_elements(1611) <= cp_elements(1229);
    -- CP-element group 1612 transition  output  bypass 
    -- predecessors 1607 
    -- successors 1613 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Sample/rr
      -- 
    cp_elements(1612) <= cp_elements(1607);
    rr_6959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1612), ack => binary_1447_inst_req_0); -- 
    -- CP-element group 1613 transition  input  no-bypass 
    -- predecessors 1612 
    -- successors 1608 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Sample/ra
      -- 
    ra_6960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1447_inst_ack_0, ack => cp_elements(1613)); -- 
    -- CP-element group 1614 transition  output  bypass 
    -- predecessors 1608 
    -- successors 1615 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Update/cr
      -- 
    cp_elements(1614) <= cp_elements(1608);
    cr_6964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1614), ack => binary_1447_inst_req_1); -- 
    -- CP-element group 1615 transition  input  no-bypass 
    -- predecessors 1614 
    -- successors 1609 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1447_complete_Update/ca
      -- 
    ca_6965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1447_inst_ack_1, ack => cp_elements(1615)); -- 
    -- CP-element group 1616 join  fork  transition  bypass 
    -- predecessors 1600 1609 
    -- successors 1617 1619 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_trigger_
      -- 
    cpelement_group_1616 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1600);
      predecessors(1) <= cp_elements(1609);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1616)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1616),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1617 join  fork  transition  no-bypass 
    -- predecessors 1616 1620 
    -- successors 1618 1621 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_active_
      -- 
    cpelement_group_1617 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1616);
      predecessors(1) <= cp_elements(1620);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1617)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1617),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1618 join  transition  no-bypass 
    -- predecessors 1617 1622 
    -- successors 1648 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1453_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1453_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1453_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1470_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1470_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1470_completed_
      -- 
    cpelement_group_1618 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1617);
      predecessors(1) <= cp_elements(1622);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1618)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1618),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1619 transition  output  bypass 
    -- predecessors 1616 
    -- successors 1620 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Sample/rr
      -- 
    cp_elements(1619) <= cp_elements(1616);
    rr_6981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1619), ack => binary_1452_inst_req_0); -- 
    -- CP-element group 1620 transition  input  no-bypass 
    -- predecessors 1619 
    -- successors 1617 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Sample/ra
      -- 
    ra_6982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1452_inst_ack_0, ack => cp_elements(1620)); -- 
    -- CP-element group 1621 transition  output  bypass 
    -- predecessors 1617 
    -- successors 1622 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Update/cr
      -- 
    cp_elements(1621) <= cp_elements(1617);
    cr_6986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1621), ack => binary_1452_inst_req_1); -- 
    -- CP-element group 1622 transition  input  no-bypass 
    -- predecessors 1621 
    -- successors 1618 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1452_complete_Update/ca
      -- 
    ca_6987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1452_inst_ack_1, ack => cp_elements(1622)); -- 
    -- CP-element group 1623 join  fork  transition  no-bypass 
    -- predecessors 1626 1627 
    -- successors 1624 1628 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_trigger_
      -- 
    cpelement_group_1623 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1626);
      predecessors(1) <= cp_elements(1627);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1623)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1623),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1624 join  fork  transition  no-bypass 
    -- predecessors 1623 1629 
    -- successors 1625 1630 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_active_
      -- 
    cpelement_group_1624 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1623);
      predecessors(1) <= cp_elements(1629);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1624)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1624),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1625 join  transition  bypass 
    -- predecessors 1624 1631 
    -- successors 1641 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1458_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1458_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1458_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1465_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1465_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1465_completed_
      -- 
    cpelement_group_1625 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1624);
      predecessors(1) <= cp_elements(1631);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1625)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1625),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1626 transition  bypass 
    -- predecessors 1449 
    -- successors 1623 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1455_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1455_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1455_completed_
      -- 
    cp_elements(1626) <= cp_elements(1449);
    -- CP-element group 1627 transition  bypass 
    -- predecessors 1239 
    -- successors 1623 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1456_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1456_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1456_completed_
      -- 
    cp_elements(1627) <= cp_elements(1239);
    -- CP-element group 1628 transition  output  bypass 
    -- predecessors 1623 
    -- successors 1629 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Sample/rr
      -- 
    cp_elements(1628) <= cp_elements(1623);
    rr_7003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1628), ack => binary_1457_inst_req_0); -- 
    -- CP-element group 1629 transition  input  no-bypass 
    -- predecessors 1628 
    -- successors 1624 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Sample/ra
      -- 
    ra_7004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1457_inst_ack_0, ack => cp_elements(1629)); -- 
    -- CP-element group 1630 transition  output  bypass 
    -- predecessors 1624 
    -- successors 1631 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Update/cr
      -- 
    cp_elements(1630) <= cp_elements(1624);
    cr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1630), ack => binary_1457_inst_req_1); -- 
    -- CP-element group 1631 transition  input  no-bypass 
    -- predecessors 1630 
    -- successors 1625 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1457_complete_Update/ca
      -- 
    ca_7009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1457_inst_ack_1, ack => cp_elements(1631)); -- 
    -- CP-element group 1632 join  fork  transition  no-bypass 
    -- predecessors 1635 1636 
    -- successors 1633 1637 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_trigger_
      -- 
    cpelement_group_1632 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1635);
      predecessors(1) <= cp_elements(1636);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1632)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1632),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1633 join  fork  transition  no-bypass 
    -- predecessors 1632 1638 
    -- successors 1634 1639 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_active_
      -- 
    cpelement_group_1633 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1632);
      predecessors(1) <= cp_elements(1638);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1633)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1633),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1634 join  transition  bypass 
    -- predecessors 1633 1640 
    -- successors 1641 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1463_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1463_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1463_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1466_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1466_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1466_completed_
      -- 
    cpelement_group_1634 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1633);
      predecessors(1) <= cp_elements(1640);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1634)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1634),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1635 transition  bypass 
    -- predecessors 1459 
    -- successors 1632 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1460_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1460_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1460_completed_
      -- 
    cp_elements(1635) <= cp_elements(1459);
    -- CP-element group 1636 transition  bypass 
    -- predecessors 1249 
    -- successors 1632 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1461_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1461_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1461_completed_
      -- 
    cp_elements(1636) <= cp_elements(1249);
    -- CP-element group 1637 transition  output  bypass 
    -- predecessors 1632 
    -- successors 1638 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Sample/rr
      -- 
    cp_elements(1637) <= cp_elements(1632);
    rr_7025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1637), ack => binary_1462_inst_req_0); -- 
    -- CP-element group 1638 transition  input  no-bypass 
    -- predecessors 1637 
    -- successors 1633 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Sample/ra
      -- 
    ra_7026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1462_inst_ack_0, ack => cp_elements(1638)); -- 
    -- CP-element group 1639 transition  output  bypass 
    -- predecessors 1633 
    -- successors 1640 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Update/cr
      -- 
    cp_elements(1639) <= cp_elements(1633);
    cr_7030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1639), ack => binary_1462_inst_req_1); -- 
    -- CP-element group 1640 transition  input  no-bypass 
    -- predecessors 1639 
    -- successors 1634 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1462_complete_Update/ca
      -- 
    ca_7031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1462_inst_ack_1, ack => cp_elements(1640)); -- 
    -- CP-element group 1641 join  fork  transition  bypass 
    -- predecessors 1625 1634 
    -- successors 1642 1644 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_trigger_
      -- 
    cpelement_group_1641 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1625);
      predecessors(1) <= cp_elements(1634);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1641)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1641),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1642 join  fork  transition  no-bypass 
    -- predecessors 1641 1645 
    -- successors 1643 1646 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_active_
      -- 
    cpelement_group_1642 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1641);
      predecessors(1) <= cp_elements(1645);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1642)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1642),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1643 join  transition  no-bypass 
    -- predecessors 1642 1647 
    -- successors 1648 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1468_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1468_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1468_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1471_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1471_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1471_completed_
      -- 
    cpelement_group_1643 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1642);
      predecessors(1) <= cp_elements(1647);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1643)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1643),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1644 transition  output  bypass 
    -- predecessors 1641 
    -- successors 1645 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Sample/rr
      -- 
    cp_elements(1644) <= cp_elements(1641);
    rr_7047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1644), ack => binary_1467_inst_req_0); -- 
    -- CP-element group 1645 transition  input  no-bypass 
    -- predecessors 1644 
    -- successors 1642 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Sample/ra
      -- 
    ra_7048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1467_inst_ack_0, ack => cp_elements(1645)); -- 
    -- CP-element group 1646 transition  output  bypass 
    -- predecessors 1642 
    -- successors 1647 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Update/cr
      -- 
    cp_elements(1646) <= cp_elements(1642);
    cr_7052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1646), ack => binary_1467_inst_req_1); -- 
    -- CP-element group 1647 transition  input  no-bypass 
    -- predecessors 1646 
    -- successors 1643 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1467_complete_Update/ca
      -- 
    ca_7053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1467_inst_ack_1, ack => cp_elements(1647)); -- 
    -- CP-element group 1648 join  fork  transition  bypass 
    -- predecessors 1618 1643 
    -- successors 1649 1651 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_trigger_
      -- 
    cpelement_group_1648 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1618);
      predecessors(1) <= cp_elements(1643);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1648)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1648),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1649 join  fork  transition  no-bypass 
    -- predecessors 1648 1652 
    -- successors 1650 1653 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_active_
      -- 
    cpelement_group_1649 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1648);
      predecessors(1) <= cp_elements(1652);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1649)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1649),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1650 join  transition  no-bypass 
    -- predecessors 1649 1654 
    -- successors 1655 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1473_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1473_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1473_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1476_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1476_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1476_completed_
      -- 
    cpelement_group_1650 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1649);
      predecessors(1) <= cp_elements(1654);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1650)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1650),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1651 transition  output  bypass 
    -- predecessors 1648 
    -- successors 1652 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Sample/rr
      -- 
    cp_elements(1651) <= cp_elements(1648);
    rr_7069_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1651), ack => binary_1472_inst_req_0); -- 
    -- CP-element group 1652 transition  input  no-bypass 
    -- predecessors 1651 
    -- successors 1649 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Sample/ra
      -- 
    ra_7070_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1472_inst_ack_0, ack => cp_elements(1652)); -- 
    -- CP-element group 1653 transition  output  bypass 
    -- predecessors 1649 
    -- successors 1654 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Update/cr
      -- 
    cp_elements(1653) <= cp_elements(1649);
    cr_7074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1653), ack => binary_1472_inst_req_1); -- 
    -- CP-element group 1654 transition  input  no-bypass 
    -- predecessors 1653 
    -- successors 1650 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1472_complete_Update/ca
      -- 
    ca_7075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1472_inst_ack_1, ack => cp_elements(1654)); -- 
    -- CP-element group 1655 join  fork  transition  no-bypass 
    -- predecessors 1650 1658 
    -- successors 1656 1659 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_trigger_
      -- 
    cpelement_group_1655 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1650);
      predecessors(1) <= cp_elements(1658);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1655)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1655),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1656 join  fork  transition  bypass 
    -- predecessors 1655 1660 
    -- successors 1657 1661 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_active_
      -- 
    cpelement_group_1656 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1655);
      predecessors(1) <= cp_elements(1660);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1656)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1656),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1657 join  transition  bypass 
    -- predecessors 1656 1662 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1478_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1478_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1478_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_completed_
      -- 
    cpelement_group_1657 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1656);
      predecessors(1) <= cp_elements(1662);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1657)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1657),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1658 transition  bypass 
    -- predecessors 367 
    -- successors 1655 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1475_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1475_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1475_completed_
      -- 
    cp_elements(1658) <= cp_elements(367);
    -- CP-element group 1659 transition  output  bypass 
    -- predecessors 1655 
    -- successors 1660 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Sample/rr
      -- 
    cp_elements(1659) <= cp_elements(1655);
    rr_7091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1659), ack => binary_1477_inst_req_0); -- 
    -- CP-element group 1660 transition  input  no-bypass 
    -- predecessors 1659 
    -- successors 1656 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Sample/ra
      -- 
    ra_7092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1477_inst_ack_0, ack => cp_elements(1660)); -- 
    -- CP-element group 1661 transition  output  bypass 
    -- predecessors 1656 
    -- successors 1662 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Update/cr
      -- 
    cp_elements(1661) <= cp_elements(1656);
    cr_7096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1661), ack => binary_1477_inst_req_1); -- 
    -- CP-element group 1662 transition  input  no-bypass 
    -- predecessors 1661 
    -- successors 1657 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1477_complete_Update/ca
      -- 
    ca_7097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1477_inst_ack_1, ack => cp_elements(1662)); -- 
    -- CP-element group 1663 join  fork  transition  no-bypass 
    -- predecessors 1666 1667 
    -- successors 1664 1668 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_trigger_
      -- 
    cpelement_group_1663 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1666);
      predecessors(1) <= cp_elements(1667);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1663)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1663),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1664 join  fork  transition  no-bypass 
    -- predecessors 1663 1669 
    -- successors 1665 1670 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_active_
      -- 
    cpelement_group_1664 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1663);
      predecessors(1) <= cp_elements(1669);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1664)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1664),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1665 join  transition  bypass 
    -- predecessors 1664 1671 
    -- successors 1681 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1483_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1483_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1483_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1490_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1490_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1490_completed_
      -- 
    cpelement_group_1665 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1664);
      predecessors(1) <= cp_elements(1671);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1665)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1665),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1666 transition  bypass 
    -- predecessors 1429 
    -- successors 1663 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1480_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1480_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1480_completed_
      -- 
    cp_elements(1666) <= cp_elements(1429);
    -- CP-element group 1667 transition  bypass 
    -- predecessors 1324 
    -- successors 1663 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1481_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1481_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1481_completed_
      -- 
    cp_elements(1667) <= cp_elements(1324);
    -- CP-element group 1668 transition  output  bypass 
    -- predecessors 1663 
    -- successors 1669 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Sample/rr
      -- 
    cp_elements(1668) <= cp_elements(1663);
    rr_7113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1668), ack => binary_1482_inst_req_0); -- 
    -- CP-element group 1669 transition  input  no-bypass 
    -- predecessors 1668 
    -- successors 1664 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Sample/ra
      -- 
    ra_7114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1482_inst_ack_0, ack => cp_elements(1669)); -- 
    -- CP-element group 1670 transition  output  bypass 
    -- predecessors 1664 
    -- successors 1671 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Update/cr
      -- 
    cp_elements(1670) <= cp_elements(1664);
    cr_7118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1670), ack => binary_1482_inst_req_1); -- 
    -- CP-element group 1671 transition  input  no-bypass 
    -- predecessors 1670 
    -- successors 1665 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1482_complete_Update/ca
      -- 
    ca_7119_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1482_inst_ack_1, ack => cp_elements(1671)); -- 
    -- CP-element group 1672 join  fork  transition  no-bypass 
    -- predecessors 1675 1676 
    -- successors 1673 1677 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_trigger_
      -- 
    cpelement_group_1672 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1675);
      predecessors(1) <= cp_elements(1676);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1672)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1672),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1673 join  fork  transition  no-bypass 
    -- predecessors 1672 1678 
    -- successors 1674 1679 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_active_
      -- 
    cpelement_group_1673 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1672);
      predecessors(1) <= cp_elements(1678);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1673)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1673),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1674 join  transition  bypass 
    -- predecessors 1673 1680 
    -- successors 1681 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1488_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1488_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1488_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1491_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1491_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1491_completed_
      -- 
    cpelement_group_1674 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1673);
      predecessors(1) <= cp_elements(1680);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1674)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1674),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1675 transition  bypass 
    -- predecessors 1439 
    -- successors 1672 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1485_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1485_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1485_completed_
      -- 
    cp_elements(1675) <= cp_elements(1439);
    -- CP-element group 1676 transition  bypass 
    -- predecessors 1334 
    -- successors 1672 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1486_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1486_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1486_completed_
      -- 
    cp_elements(1676) <= cp_elements(1334);
    -- CP-element group 1677 transition  output  bypass 
    -- predecessors 1672 
    -- successors 1678 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Sample/rr
      -- 
    cp_elements(1677) <= cp_elements(1672);
    rr_7135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1677), ack => binary_1487_inst_req_0); -- 
    -- CP-element group 1678 transition  input  no-bypass 
    -- predecessors 1677 
    -- successors 1673 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Sample/ra
      -- 
    ra_7136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1487_inst_ack_0, ack => cp_elements(1678)); -- 
    -- CP-element group 1679 transition  output  bypass 
    -- predecessors 1673 
    -- successors 1680 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Update/cr
      -- 
    cp_elements(1679) <= cp_elements(1673);
    cr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1679), ack => binary_1487_inst_req_1); -- 
    -- CP-element group 1680 transition  input  no-bypass 
    -- predecessors 1679 
    -- successors 1674 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1487_complete_Update/ca
      -- 
    ca_7141_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1487_inst_ack_1, ack => cp_elements(1680)); -- 
    -- CP-element group 1681 join  fork  transition  bypass 
    -- predecessors 1665 1674 
    -- successors 1682 1684 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_trigger_
      -- 
    cpelement_group_1681 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1665);
      predecessors(1) <= cp_elements(1674);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1681)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1681),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1682 join  fork  transition  no-bypass 
    -- predecessors 1681 1685 
    -- successors 1683 1686 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_active_
      -- 
    cpelement_group_1682 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1681);
      predecessors(1) <= cp_elements(1685);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1682)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1682),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1683 join  transition  no-bypass 
    -- predecessors 1682 1687 
    -- successors 1713 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1493_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1493_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1493_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1510_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1510_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1510_completed_
      -- 
    cpelement_group_1683 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1682);
      predecessors(1) <= cp_elements(1687);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1683)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1683),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1684 transition  output  bypass 
    -- predecessors 1681 
    -- successors 1685 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Sample/rr
      -- 
    cp_elements(1684) <= cp_elements(1681);
    rr_7157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1684), ack => binary_1492_inst_req_0); -- 
    -- CP-element group 1685 transition  input  no-bypass 
    -- predecessors 1684 
    -- successors 1682 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Sample/ra
      -- 
    ra_7158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1492_inst_ack_0, ack => cp_elements(1685)); -- 
    -- CP-element group 1686 transition  output  bypass 
    -- predecessors 1682 
    -- successors 1687 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Update/cr
      -- 
    cp_elements(1686) <= cp_elements(1682);
    cr_7162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1686), ack => binary_1492_inst_req_1); -- 
    -- CP-element group 1687 transition  input  no-bypass 
    -- predecessors 1686 
    -- successors 1683 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1492_complete_Update/ca
      -- 
    ca_7163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1492_inst_ack_1, ack => cp_elements(1687)); -- 
    -- CP-element group 1688 join  fork  transition  no-bypass 
    -- predecessors 1691 1692 
    -- successors 1689 1693 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_trigger_
      -- 
    cpelement_group_1688 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1691);
      predecessors(1) <= cp_elements(1692);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1688)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1688),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1689 join  fork  transition  no-bypass 
    -- predecessors 1688 1694 
    -- successors 1690 1695 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_active_
      -- 
    cpelement_group_1689 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1688);
      predecessors(1) <= cp_elements(1694);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1689)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1689),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1690 join  transition  bypass 
    -- predecessors 1689 1696 
    -- successors 1706 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1498_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1498_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1498_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1505_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1505_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1505_completed_
      -- 
    cpelement_group_1690 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1689);
      predecessors(1) <= cp_elements(1696);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1690)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1690),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1691 transition  bypass 
    -- predecessors 1449 
    -- successors 1688 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1495_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1495_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1495_completed_
      -- 
    cp_elements(1691) <= cp_elements(1449);
    -- CP-element group 1692 transition  bypass 
    -- predecessors 1344 
    -- successors 1688 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1496_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1496_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1496_completed_
      -- 
    cp_elements(1692) <= cp_elements(1344);
    -- CP-element group 1693 transition  output  bypass 
    -- predecessors 1688 
    -- successors 1694 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Sample/rr
      -- 
    cp_elements(1693) <= cp_elements(1688);
    rr_7179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1693), ack => binary_1497_inst_req_0); -- 
    -- CP-element group 1694 transition  input  no-bypass 
    -- predecessors 1693 
    -- successors 1689 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Sample/ra
      -- 
    ra_7180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1497_inst_ack_0, ack => cp_elements(1694)); -- 
    -- CP-element group 1695 transition  output  bypass 
    -- predecessors 1689 
    -- successors 1696 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Update/cr
      -- 
    cp_elements(1695) <= cp_elements(1689);
    cr_7184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1695), ack => binary_1497_inst_req_1); -- 
    -- CP-element group 1696 transition  input  no-bypass 
    -- predecessors 1695 
    -- successors 1690 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1497_complete_Update/ca
      -- 
    ca_7185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1497_inst_ack_1, ack => cp_elements(1696)); -- 
    -- CP-element group 1697 join  fork  transition  no-bypass 
    -- predecessors 1700 1701 
    -- successors 1698 1702 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_trigger_
      -- 
    cpelement_group_1697 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1700);
      predecessors(1) <= cp_elements(1701);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1697)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1697),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1698 join  fork  transition  no-bypass 
    -- predecessors 1697 1703 
    -- successors 1699 1704 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_active_
      -- 
    cpelement_group_1698 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1697);
      predecessors(1) <= cp_elements(1703);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1698)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1698),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1699 join  transition  bypass 
    -- predecessors 1698 1705 
    -- successors 1706 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1503_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1503_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1503_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1506_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1506_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1506_completed_
      -- 
    cpelement_group_1699 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1698);
      predecessors(1) <= cp_elements(1705);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1699)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1699),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1700 transition  bypass 
    -- predecessors 1459 
    -- successors 1697 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1500_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1500_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1500_completed_
      -- 
    cp_elements(1700) <= cp_elements(1459);
    -- CP-element group 1701 transition  bypass 
    -- predecessors 1354 
    -- successors 1697 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1501_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1501_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1501_completed_
      -- 
    cp_elements(1701) <= cp_elements(1354);
    -- CP-element group 1702 transition  output  bypass 
    -- predecessors 1697 
    -- successors 1703 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Sample/rr
      -- 
    cp_elements(1702) <= cp_elements(1697);
    rr_7201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1702), ack => binary_1502_inst_req_0); -- 
    -- CP-element group 1703 transition  input  no-bypass 
    -- predecessors 1702 
    -- successors 1698 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Sample/ra
      -- 
    ra_7202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1502_inst_ack_0, ack => cp_elements(1703)); -- 
    -- CP-element group 1704 transition  output  bypass 
    -- predecessors 1698 
    -- successors 1705 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Update/cr
      -- 
    cp_elements(1704) <= cp_elements(1698);
    cr_7206_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1704), ack => binary_1502_inst_req_1); -- 
    -- CP-element group 1705 transition  input  no-bypass 
    -- predecessors 1704 
    -- successors 1699 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1502_complete_Update/ca
      -- 
    ca_7207_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1502_inst_ack_1, ack => cp_elements(1705)); -- 
    -- CP-element group 1706 join  fork  transition  bypass 
    -- predecessors 1690 1699 
    -- successors 1707 1709 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_trigger_
      -- 
    cpelement_group_1706 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1690);
      predecessors(1) <= cp_elements(1699);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1706)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1706),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1707 join  fork  transition  no-bypass 
    -- predecessors 1706 1710 
    -- successors 1708 1711 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_active_
      -- 
    cpelement_group_1707 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1706);
      predecessors(1) <= cp_elements(1710);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1707)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1707),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1708 join  transition  no-bypass 
    -- predecessors 1707 1712 
    -- successors 1713 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1508_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1508_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1508_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1511_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1511_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1511_completed_
      -- 
    cpelement_group_1708 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1707);
      predecessors(1) <= cp_elements(1712);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1708)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1708),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1709 transition  output  bypass 
    -- predecessors 1706 
    -- successors 1710 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Sample/rr
      -- 
    cp_elements(1709) <= cp_elements(1706);
    rr_7223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1709), ack => binary_1507_inst_req_0); -- 
    -- CP-element group 1710 transition  input  no-bypass 
    -- predecessors 1709 
    -- successors 1707 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Sample/ra
      -- 
    ra_7224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1507_inst_ack_0, ack => cp_elements(1710)); -- 
    -- CP-element group 1711 transition  output  bypass 
    -- predecessors 1707 
    -- successors 1712 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Update/cr
      -- 
    cp_elements(1711) <= cp_elements(1707);
    cr_7228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1711), ack => binary_1507_inst_req_1); -- 
    -- CP-element group 1712 transition  input  no-bypass 
    -- predecessors 1711 
    -- successors 1708 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1507_complete_Update/ca
      -- 
    ca_7229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1507_inst_ack_1, ack => cp_elements(1712)); -- 
    -- CP-element group 1713 join  fork  transition  bypass 
    -- predecessors 1683 1708 
    -- successors 1714 1716 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_trigger_
      -- 
    cpelement_group_1713 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1683);
      predecessors(1) <= cp_elements(1708);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1713)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1713),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1714 join  fork  transition  no-bypass 
    -- predecessors 1713 1717 
    -- successors 1715 1718 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_active_
      -- 
    cpelement_group_1714 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1713);
      predecessors(1) <= cp_elements(1717);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1714)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1714),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1715 join  transition  no-bypass 
    -- predecessors 1714 1719 
    -- successors 1720 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1513_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1513_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1513_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1516_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1516_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1516_completed_
      -- 
    cpelement_group_1715 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1714);
      predecessors(1) <= cp_elements(1719);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1715)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1715),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1716 transition  output  bypass 
    -- predecessors 1713 
    -- successors 1717 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Sample/rr
      -- 
    cp_elements(1716) <= cp_elements(1713);
    rr_7245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1716), ack => binary_1512_inst_req_0); -- 
    -- CP-element group 1717 transition  input  no-bypass 
    -- predecessors 1716 
    -- successors 1714 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Sample/ra
      -- 
    ra_7246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1512_inst_ack_0, ack => cp_elements(1717)); -- 
    -- CP-element group 1718 transition  output  bypass 
    -- predecessors 1714 
    -- successors 1719 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Update/cr
      -- 
    cp_elements(1718) <= cp_elements(1714);
    cr_7250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1718), ack => binary_1512_inst_req_1); -- 
    -- CP-element group 1719 transition  input  no-bypass 
    -- predecessors 1718 
    -- successors 1715 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1512_complete_Update/ca
      -- 
    ca_7251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1512_inst_ack_1, ack => cp_elements(1719)); -- 
    -- CP-element group 1720 join  fork  transition  no-bypass 
    -- predecessors 1715 1723 
    -- successors 1721 1724 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_trigger_
      -- 
    cpelement_group_1720 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1715);
      predecessors(1) <= cp_elements(1723);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1720)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1720),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1721 join  fork  transition  bypass 
    -- predecessors 1720 1725 
    -- successors 1722 1726 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_active_
      -- 
    cpelement_group_1721 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1720);
      predecessors(1) <= cp_elements(1725);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1721)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1721),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1722 join  transition  bypass 
    -- predecessors 1721 1727 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1518_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1518_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1518_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_completed_
      -- 
    cpelement_group_1722 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1721);
      predecessors(1) <= cp_elements(1727);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1722)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1722),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1723 transition  bypass 
    -- predecessors 367 
    -- successors 1720 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1515_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1515_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1515_completed_
      -- 
    cp_elements(1723) <= cp_elements(367);
    -- CP-element group 1724 transition  output  bypass 
    -- predecessors 1720 
    -- successors 1725 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Sample/rr
      -- 
    cp_elements(1724) <= cp_elements(1720);
    rr_7267_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1724), ack => binary_1517_inst_req_0); -- 
    -- CP-element group 1725 transition  input  no-bypass 
    -- predecessors 1724 
    -- successors 1721 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Sample/ra
      -- 
    ra_7268_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1517_inst_ack_0, ack => cp_elements(1725)); -- 
    -- CP-element group 1726 transition  output  bypass 
    -- predecessors 1721 
    -- successors 1727 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Update/cr
      -- 
    cp_elements(1726) <= cp_elements(1721);
    cr_7272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1726), ack => binary_1517_inst_req_1); -- 
    -- CP-element group 1727 transition  input  no-bypass 
    -- predecessors 1726 
    -- successors 1722 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1517_complete_Update/ca
      -- 
    ca_7273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1517_inst_ack_1, ack => cp_elements(1727)); -- 
    -- CP-element group 1728 join  fork  transition  bypass 
    -- predecessors 1732 1734 
    -- successors 1729 1735 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_active_
      -- 
    cpelement_group_1728 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1732);
      predecessors(1) <= cp_elements(1734);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1728)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1728),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1729 join  fork  transition  bypass 
    -- predecessors 1728 1737 
    -- successors 1771 1836 1901 1966 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1522_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1522_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1522_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_completed_
      -- 
    cpelement_group_1729 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1728);
      predecessors(1) <= cp_elements(1737);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1729)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1729),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1730 transition  input  output  no-bypass 
    -- predecessors 517 
    -- successors 1731 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7291_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1521_base_resize_ack_0, ack => cp_elements(1730)); -- 
    sum_rename_req_7295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1730), ack => ptr_deref_1521_root_address_inst_req_0); -- 
    -- CP-element group 1731 transition  input  output  no-bypass 
    -- predecessors 1730 
    -- successors 1732 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1521_root_address_inst_ack_0, ack => cp_elements(1731)); -- 
    root_register_req_7300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1731), ack => ptr_deref_1521_addr_0_req_0); -- 
    -- CP-element group 1732 fork  transition  input  no-bypass 
    -- predecessors 1731 
    -- successors 1728 1733 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_word_addrgen/root_register_ack
      -- 
    root_register_ack_7301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1521_addr_0_ack_0, ack => cp_elements(1732)); -- 
    -- CP-element group 1733 transition  output  bypass 
    -- predecessors 1732 
    -- successors 1734 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/word_access/word_access_0/rr
      -- 
    cp_elements(1733) <= cp_elements(1732);
    rr_7311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1733), ack => ptr_deref_1521_load_0_req_0); -- 
    -- CP-element group 1734 transition  input  no-bypass 
    -- predecessors 1733 
    -- successors 1728 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_request/word_access/word_access_0/ra
      -- 
    ra_7312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1521_load_0_ack_0, ack => cp_elements(1734)); -- 
    -- CP-element group 1735 transition  output  bypass 
    -- predecessors 1728 
    -- successors 1736 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1735) <= cp_elements(1728);
    cr_7322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1735), ack => ptr_deref_1521_load_0_req_1); -- 
    -- CP-element group 1736 transition  input  output  no-bypass 
    -- predecessors 1735 
    -- successors 1737 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/merge_req
      -- 
    ca_7323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1521_load_0_ack_1, ack => cp_elements(1736)); -- 
    merge_req_7324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1736), ack => ptr_deref_1521_gather_scatter_req_0); -- 
    -- CP-element group 1737 transition  input  no-bypass 
    -- predecessors 1736 
    -- successors 1729 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1521_complete/merge_ack
      -- 
    merge_ack_7325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1521_gather_scatter_ack_0, ack => cp_elements(1737)); -- 
    -- CP-element group 1738 join  fork  transition  bypass 
    -- predecessors 1742 1744 
    -- successors 1739 1745 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_active_
      -- 
    cpelement_group_1738 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1742);
      predecessors(1) <= cp_elements(1744);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1738)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1738),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1739 join  fork  transition  bypass 
    -- predecessors 1738 1747 
    -- successors 1780 1845 1910 1975 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1526_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1526_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1526_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_completed_
      -- 
    cpelement_group_1739 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1738);
      predecessors(1) <= cp_elements(1747);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1739)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1739),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1740 transition  input  output  no-bypass 
    -- predecessors 568 
    -- successors 1741 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1525_base_resize_ack_0, ack => cp_elements(1740)); -- 
    sum_rename_req_7347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1740), ack => ptr_deref_1525_root_address_inst_req_0); -- 
    -- CP-element group 1741 transition  input  output  no-bypass 
    -- predecessors 1740 
    -- successors 1742 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1525_root_address_inst_ack_0, ack => cp_elements(1741)); -- 
    root_register_req_7352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1741), ack => ptr_deref_1525_addr_0_req_0); -- 
    -- CP-element group 1742 fork  transition  input  no-bypass 
    -- predecessors 1741 
    -- successors 1738 1743 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_word_addrgen/root_register_ack
      -- 
    root_register_ack_7353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1525_addr_0_ack_0, ack => cp_elements(1742)); -- 
    -- CP-element group 1743 transition  output  bypass 
    -- predecessors 1742 
    -- successors 1744 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/word_access/word_access_0/rr
      -- 
    cp_elements(1743) <= cp_elements(1742);
    rr_7363_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1743), ack => ptr_deref_1525_load_0_req_0); -- 
    -- CP-element group 1744 transition  input  no-bypass 
    -- predecessors 1743 
    -- successors 1738 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_request/word_access/word_access_0/ra
      -- 
    ra_7364_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1525_load_0_ack_0, ack => cp_elements(1744)); -- 
    -- CP-element group 1745 transition  output  bypass 
    -- predecessors 1738 
    -- successors 1746 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1745) <= cp_elements(1738);
    cr_7374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1745), ack => ptr_deref_1525_load_0_req_1); -- 
    -- CP-element group 1746 transition  input  output  no-bypass 
    -- predecessors 1745 
    -- successors 1747 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/merge_req
      -- 
    ca_7375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1525_load_0_ack_1, ack => cp_elements(1746)); -- 
    merge_req_7376_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1746), ack => ptr_deref_1525_gather_scatter_req_0); -- 
    -- CP-element group 1747 transition  input  no-bypass 
    -- predecessors 1746 
    -- successors 1739 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1525_complete/merge_ack
      -- 
    merge_ack_7377_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1525_gather_scatter_ack_0, ack => cp_elements(1747)); -- 
    -- CP-element group 1748 join  fork  transition  bypass 
    -- predecessors 1752 1754 
    -- successors 1749 1755 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_active_
      -- 
    cpelement_group_1748 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1752);
      predecessors(1) <= cp_elements(1754);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1748)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1748),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1749 join  fork  transition  bypass 
    -- predecessors 1748 1757 
    -- successors 1796 1861 1926 1991 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1530_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1530_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1530_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_completed_
      -- 
    cpelement_group_1749 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1748);
      predecessors(1) <= cp_elements(1757);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1749)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1749),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1750 transition  input  output  no-bypass 
    -- predecessors 551 
    -- successors 1751 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7395_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_base_resize_ack_0, ack => cp_elements(1750)); -- 
    sum_rename_req_7399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1750), ack => ptr_deref_1529_root_address_inst_req_0); -- 
    -- CP-element group 1751 transition  input  output  no-bypass 
    -- predecessors 1750 
    -- successors 1752 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_root_address_inst_ack_0, ack => cp_elements(1751)); -- 
    root_register_req_7404_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1751), ack => ptr_deref_1529_addr_0_req_0); -- 
    -- CP-element group 1752 fork  transition  input  no-bypass 
    -- predecessors 1751 
    -- successors 1748 1753 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_word_addrgen/root_register_ack
      -- 
    root_register_ack_7405_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_addr_0_ack_0, ack => cp_elements(1752)); -- 
    -- CP-element group 1753 transition  output  bypass 
    -- predecessors 1752 
    -- successors 1754 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/word_access/word_access_0/rr
      -- 
    cp_elements(1753) <= cp_elements(1752);
    rr_7415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1753), ack => ptr_deref_1529_load_0_req_0); -- 
    -- CP-element group 1754 transition  input  no-bypass 
    -- predecessors 1753 
    -- successors 1748 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_request/word_access/word_access_0/ra
      -- 
    ra_7416_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_load_0_ack_0, ack => cp_elements(1754)); -- 
    -- CP-element group 1755 transition  output  bypass 
    -- predecessors 1748 
    -- successors 1756 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1755) <= cp_elements(1748);
    cr_7426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1755), ack => ptr_deref_1529_load_0_req_1); -- 
    -- CP-element group 1756 transition  input  output  no-bypass 
    -- predecessors 1755 
    -- successors 1757 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/merge_req
      -- 
    ca_7427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_load_0_ack_1, ack => cp_elements(1756)); -- 
    merge_req_7428_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1756), ack => ptr_deref_1529_gather_scatter_req_0); -- 
    -- CP-element group 1757 transition  input  no-bypass 
    -- predecessors 1756 
    -- successors 1749 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1529_complete/merge_ack
      -- 
    merge_ack_7429_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_gather_scatter_ack_0, ack => cp_elements(1757)); -- 
    -- CP-element group 1758 join  fork  transition  bypass 
    -- predecessors 1762 1764 
    -- successors 1759 1765 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_active_
      -- 
    cpelement_group_1758 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1762);
      predecessors(1) <= cp_elements(1764);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1758)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1758),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1759 join  fork  transition  bypass 
    -- predecessors 1758 1767 
    -- successors 1805 1870 1935 2000 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1534_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1534_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1534_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_completed_
      -- 
    cpelement_group_1759 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1758);
      predecessors(1) <= cp_elements(1767);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1759)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1759),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1760 transition  input  output  no-bypass 
    -- predecessors 534 
    -- successors 1761 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7447_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_base_resize_ack_0, ack => cp_elements(1760)); -- 
    sum_rename_req_7451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1760), ack => ptr_deref_1533_root_address_inst_req_0); -- 
    -- CP-element group 1761 transition  input  output  no-bypass 
    -- predecessors 1760 
    -- successors 1762 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_root_address_inst_ack_0, ack => cp_elements(1761)); -- 
    root_register_req_7456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1761), ack => ptr_deref_1533_addr_0_req_0); -- 
    -- CP-element group 1762 fork  transition  input  no-bypass 
    -- predecessors 1761 
    -- successors 1758 1763 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_word_addrgen/root_register_ack
      -- 
    root_register_ack_7457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_addr_0_ack_0, ack => cp_elements(1762)); -- 
    -- CP-element group 1763 transition  output  bypass 
    -- predecessors 1762 
    -- successors 1764 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/word_access/word_access_0/rr
      -- 
    cp_elements(1763) <= cp_elements(1762);
    rr_7467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1763), ack => ptr_deref_1533_load_0_req_0); -- 
    -- CP-element group 1764 transition  input  no-bypass 
    -- predecessors 1763 
    -- successors 1758 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_request/word_access/word_access_0/ra
      -- 
    ra_7468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_load_0_ack_0, ack => cp_elements(1764)); -- 
    -- CP-element group 1765 transition  output  bypass 
    -- predecessors 1758 
    -- successors 1766 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1765) <= cp_elements(1758);
    cr_7478_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1765), ack => ptr_deref_1533_load_0_req_1); -- 
    -- CP-element group 1766 transition  input  output  no-bypass 
    -- predecessors 1765 
    -- successors 1767 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/merge_req
      -- 
    ca_7479_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_load_0_ack_1, ack => cp_elements(1766)); -- 
    merge_req_7480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1766), ack => ptr_deref_1533_gather_scatter_req_0); -- 
    -- CP-element group 1767 transition  input  no-bypass 
    -- predecessors 1766 
    -- successors 1759 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1533_complete/merge_ack
      -- 
    merge_ack_7481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1533_gather_scatter_ack_0, ack => cp_elements(1767)); -- 
    -- CP-element group 1768 join  fork  transition  no-bypass 
    -- predecessors 1771 1772 
    -- successors 1769 1773 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_trigger_
      -- 
    cpelement_group_1768 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1771);
      predecessors(1) <= cp_elements(1772);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1768)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1768),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1769 join  fork  transition  no-bypass 
    -- predecessors 1768 1774 
    -- successors 1770 1775 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_active_
      -- 
    cpelement_group_1769 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1768);
      predecessors(1) <= cp_elements(1774);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1769)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1769),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1770 join  transition  bypass 
    -- predecessors 1769 1776 
    -- successors 1786 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1539_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1539_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1539_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1546_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1546_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1546_completed_
      -- 
    cpelement_group_1770 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1769);
      predecessors(1) <= cp_elements(1776);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1770)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1770),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1771 transition  bypass 
    -- predecessors 1729 
    -- successors 1768 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1536_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1536_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1536_completed_
      -- 
    cp_elements(1771) <= cp_elements(1729);
    -- CP-element group 1772 transition  bypass 
    -- predecessors 979 
    -- successors 1768 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1537_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1537_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1537_completed_
      -- 
    cp_elements(1772) <= cp_elements(979);
    -- CP-element group 1773 transition  output  bypass 
    -- predecessors 1768 
    -- successors 1774 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Sample/rr
      -- 
    cp_elements(1773) <= cp_elements(1768);
    rr_7497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1773), ack => binary_1538_inst_req_0); -- 
    -- CP-element group 1774 transition  input  no-bypass 
    -- predecessors 1773 
    -- successors 1769 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Sample/ra
      -- 
    ra_7498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1538_inst_ack_0, ack => cp_elements(1774)); -- 
    -- CP-element group 1775 transition  output  bypass 
    -- predecessors 1769 
    -- successors 1776 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Update/cr
      -- 
    cp_elements(1775) <= cp_elements(1769);
    cr_7502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1775), ack => binary_1538_inst_req_1); -- 
    -- CP-element group 1776 transition  input  no-bypass 
    -- predecessors 1775 
    -- successors 1770 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1538_complete_Update/ca
      -- 
    ca_7503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1538_inst_ack_1, ack => cp_elements(1776)); -- 
    -- CP-element group 1777 join  fork  transition  no-bypass 
    -- predecessors 1780 1781 
    -- successors 1778 1782 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_trigger_
      -- 
    cpelement_group_1777 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1780);
      predecessors(1) <= cp_elements(1781);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1777)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1777),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1778 join  fork  transition  no-bypass 
    -- predecessors 1777 1783 
    -- successors 1779 1784 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_active_
      -- 
    cpelement_group_1778 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1777);
      predecessors(1) <= cp_elements(1783);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1778)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1778),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1779 join  transition  bypass 
    -- predecessors 1778 1785 
    -- successors 1786 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1544_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1544_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1544_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1547_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1547_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1547_completed_
      -- 
    cpelement_group_1779 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1778);
      predecessors(1) <= cp_elements(1785);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1779)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1779),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1780 transition  bypass 
    -- predecessors 1739 
    -- successors 1777 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1541_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1541_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1541_completed_
      -- 
    cp_elements(1780) <= cp_elements(1739);
    -- CP-element group 1781 transition  bypass 
    -- predecessors 999 
    -- successors 1777 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1542_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1542_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1542_completed_
      -- 
    cp_elements(1781) <= cp_elements(999);
    -- CP-element group 1782 transition  output  bypass 
    -- predecessors 1777 
    -- successors 1783 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Sample/rr
      -- 
    cp_elements(1782) <= cp_elements(1777);
    rr_7519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1782), ack => binary_1543_inst_req_0); -- 
    -- CP-element group 1783 transition  input  no-bypass 
    -- predecessors 1782 
    -- successors 1778 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Sample/ra
      -- 
    ra_7520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1543_inst_ack_0, ack => cp_elements(1783)); -- 
    -- CP-element group 1784 transition  output  bypass 
    -- predecessors 1778 
    -- successors 1785 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Update/cr
      -- 
    cp_elements(1784) <= cp_elements(1778);
    cr_7524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1784), ack => binary_1543_inst_req_1); -- 
    -- CP-element group 1785 transition  input  no-bypass 
    -- predecessors 1784 
    -- successors 1779 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1543_complete_Update/ca
      -- 
    ca_7525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1543_inst_ack_1, ack => cp_elements(1785)); -- 
    -- CP-element group 1786 join  fork  transition  bypass 
    -- predecessors 1770 1779 
    -- successors 1787 1789 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_trigger_
      -- 
    cpelement_group_1786 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1770);
      predecessors(1) <= cp_elements(1779);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1786)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1786),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1787 join  fork  transition  no-bypass 
    -- predecessors 1786 1790 
    -- successors 1788 1791 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_active_
      -- 
    cpelement_group_1787 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1786);
      predecessors(1) <= cp_elements(1790);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1787)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1787),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1788 join  transition  no-bypass 
    -- predecessors 1787 1792 
    -- successors 1818 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1549_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1549_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1549_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1566_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1566_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1566_completed_
      -- 
    cpelement_group_1788 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1787);
      predecessors(1) <= cp_elements(1792);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1788)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1788),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1789 transition  output  bypass 
    -- predecessors 1786 
    -- successors 1790 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Sample/rr
      -- 
    cp_elements(1789) <= cp_elements(1786);
    rr_7541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1789), ack => binary_1548_inst_req_0); -- 
    -- CP-element group 1790 transition  input  no-bypass 
    -- predecessors 1789 
    -- successors 1787 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Sample/ra
      -- 
    ra_7542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1548_inst_ack_0, ack => cp_elements(1790)); -- 
    -- CP-element group 1791 transition  output  bypass 
    -- predecessors 1787 
    -- successors 1792 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Update/cr
      -- 
    cp_elements(1791) <= cp_elements(1787);
    cr_7546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1791), ack => binary_1548_inst_req_1); -- 
    -- CP-element group 1792 transition  input  no-bypass 
    -- predecessors 1791 
    -- successors 1788 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1548_complete_Update/ca
      -- 
    ca_7547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1548_inst_ack_1, ack => cp_elements(1792)); -- 
    -- CP-element group 1793 join  fork  transition  no-bypass 
    -- predecessors 1796 1797 
    -- successors 1794 1798 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_trigger_
      -- 
    cpelement_group_1793 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1796);
      predecessors(1) <= cp_elements(1797);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1793)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1793),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1794 join  fork  transition  no-bypass 
    -- predecessors 1793 1799 
    -- successors 1795 1800 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_active_
      -- 
    cpelement_group_1794 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1793);
      predecessors(1) <= cp_elements(1799);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1794)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1794),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1795 join  transition  bypass 
    -- predecessors 1794 1801 
    -- successors 1811 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1554_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1554_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1554_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1561_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1561_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1561_completed_
      -- 
    cpelement_group_1795 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1794);
      predecessors(1) <= cp_elements(1801);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1795)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1795),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1796 transition  bypass 
    -- predecessors 1749 
    -- successors 1793 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1551_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1551_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1551_completed_
      -- 
    cp_elements(1796) <= cp_elements(1749);
    -- CP-element group 1797 transition  bypass 
    -- predecessors 1019 
    -- successors 1793 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1552_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1552_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1552_completed_
      -- 
    cp_elements(1797) <= cp_elements(1019);
    -- CP-element group 1798 transition  output  bypass 
    -- predecessors 1793 
    -- successors 1799 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Sample/rr
      -- 
    cp_elements(1798) <= cp_elements(1793);
    rr_7563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1798), ack => binary_1553_inst_req_0); -- 
    -- CP-element group 1799 transition  input  no-bypass 
    -- predecessors 1798 
    -- successors 1794 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Sample/ra
      -- 
    ra_7564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1553_inst_ack_0, ack => cp_elements(1799)); -- 
    -- CP-element group 1800 transition  output  bypass 
    -- predecessors 1794 
    -- successors 1801 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Update/cr
      -- 
    cp_elements(1800) <= cp_elements(1794);
    cr_7568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1800), ack => binary_1553_inst_req_1); -- 
    -- CP-element group 1801 transition  input  no-bypass 
    -- predecessors 1800 
    -- successors 1795 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1553_complete_Update/ca
      -- 
    ca_7569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1553_inst_ack_1, ack => cp_elements(1801)); -- 
    -- CP-element group 1802 join  fork  transition  no-bypass 
    -- predecessors 1805 1806 
    -- successors 1803 1807 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_trigger_
      -- 
    cpelement_group_1802 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1805);
      predecessors(1) <= cp_elements(1806);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1802)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1802),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1803 join  fork  transition  no-bypass 
    -- predecessors 1802 1808 
    -- successors 1804 1809 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_active_
      -- 
    cpelement_group_1803 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1802);
      predecessors(1) <= cp_elements(1808);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1803)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1803),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1804 join  transition  bypass 
    -- predecessors 1803 1810 
    -- successors 1811 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1559_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1559_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1559_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1562_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1562_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1562_completed_
      -- 
    cpelement_group_1804 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1803);
      predecessors(1) <= cp_elements(1810);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1804)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1804),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1805 transition  bypass 
    -- predecessors 1759 
    -- successors 1802 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1556_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1556_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1556_completed_
      -- 
    cp_elements(1805) <= cp_elements(1759);
    -- CP-element group 1806 transition  bypass 
    -- predecessors 1039 
    -- successors 1802 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1557_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1557_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1557_completed_
      -- 
    cp_elements(1806) <= cp_elements(1039);
    -- CP-element group 1807 transition  output  bypass 
    -- predecessors 1802 
    -- successors 1808 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Sample/rr
      -- 
    cp_elements(1807) <= cp_elements(1802);
    rr_7585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1807), ack => binary_1558_inst_req_0); -- 
    -- CP-element group 1808 transition  input  no-bypass 
    -- predecessors 1807 
    -- successors 1803 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Sample/ra
      -- 
    ra_7586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1558_inst_ack_0, ack => cp_elements(1808)); -- 
    -- CP-element group 1809 transition  output  bypass 
    -- predecessors 1803 
    -- successors 1810 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Update/cr
      -- 
    cp_elements(1809) <= cp_elements(1803);
    cr_7590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1809), ack => binary_1558_inst_req_1); -- 
    -- CP-element group 1810 transition  input  no-bypass 
    -- predecessors 1809 
    -- successors 1804 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1558_complete_Update/ca
      -- 
    ca_7591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1558_inst_ack_1, ack => cp_elements(1810)); -- 
    -- CP-element group 1811 join  fork  transition  bypass 
    -- predecessors 1795 1804 
    -- successors 1812 1814 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_trigger_
      -- 
    cpelement_group_1811 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1795);
      predecessors(1) <= cp_elements(1804);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1811)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1811),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1812 join  fork  transition  no-bypass 
    -- predecessors 1811 1815 
    -- successors 1813 1816 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_active_
      -- 
    cpelement_group_1812 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1811);
      predecessors(1) <= cp_elements(1815);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1812)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1812),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1813 join  transition  no-bypass 
    -- predecessors 1812 1817 
    -- successors 1818 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1564_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1564_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1564_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1567_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1567_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1567_completed_
      -- 
    cpelement_group_1813 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1812);
      predecessors(1) <= cp_elements(1817);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1813)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1813),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1814 transition  output  bypass 
    -- predecessors 1811 
    -- successors 1815 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Sample/rr
      -- 
    cp_elements(1814) <= cp_elements(1811);
    rr_7607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1814), ack => binary_1563_inst_req_0); -- 
    -- CP-element group 1815 transition  input  no-bypass 
    -- predecessors 1814 
    -- successors 1812 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Sample/ra
      -- 
    ra_7608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1563_inst_ack_0, ack => cp_elements(1815)); -- 
    -- CP-element group 1816 transition  output  bypass 
    -- predecessors 1812 
    -- successors 1817 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Update/cr
      -- 
    cp_elements(1816) <= cp_elements(1812);
    cr_7612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1816), ack => binary_1563_inst_req_1); -- 
    -- CP-element group 1817 transition  input  no-bypass 
    -- predecessors 1816 
    -- successors 1813 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1563_complete_Update/ca
      -- 
    ca_7613_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1563_inst_ack_1, ack => cp_elements(1817)); -- 
    -- CP-element group 1818 join  fork  transition  bypass 
    -- predecessors 1788 1813 
    -- successors 1819 1821 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_trigger_
      -- 
    cpelement_group_1818 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1788);
      predecessors(1) <= cp_elements(1813);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1818)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1818),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1819 join  fork  transition  no-bypass 
    -- predecessors 1818 1822 
    -- successors 1820 1823 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_active_
      -- 
    cpelement_group_1819 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1818);
      predecessors(1) <= cp_elements(1822);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1819)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1819),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1820 join  transition  no-bypass 
    -- predecessors 1819 1824 
    -- successors 1825 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1569_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1569_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1569_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1572_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1572_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1572_completed_
      -- 
    cpelement_group_1820 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1819);
      predecessors(1) <= cp_elements(1824);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1820)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1820),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1821 transition  output  bypass 
    -- predecessors 1818 
    -- successors 1822 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Sample/rr
      -- 
    cp_elements(1821) <= cp_elements(1818);
    rr_7629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1821), ack => binary_1568_inst_req_0); -- 
    -- CP-element group 1822 transition  input  no-bypass 
    -- predecessors 1821 
    -- successors 1819 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Sample/ra
      -- 
    ra_7630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1568_inst_ack_0, ack => cp_elements(1822)); -- 
    -- CP-element group 1823 transition  output  bypass 
    -- predecessors 1819 
    -- successors 1824 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Update/cr
      -- 
    cp_elements(1823) <= cp_elements(1819);
    cr_7634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1823), ack => binary_1568_inst_req_1); -- 
    -- CP-element group 1824 transition  input  no-bypass 
    -- predecessors 1823 
    -- successors 1820 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1568_complete_Update/ca
      -- 
    ca_7635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1568_inst_ack_1, ack => cp_elements(1824)); -- 
    -- CP-element group 1825 join  fork  transition  no-bypass 
    -- predecessors 1820 1828 
    -- successors 1826 1829 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_trigger_
      -- 
    cpelement_group_1825 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1820);
      predecessors(1) <= cp_elements(1828);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1825)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1825),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1826 join  fork  transition  bypass 
    -- predecessors 1825 1830 
    -- successors 1827 1831 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_active_
      -- 
    cpelement_group_1826 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1825);
      predecessors(1) <= cp_elements(1830);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1826)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1826),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1827 join  transition  bypass 
    -- predecessors 1826 1832 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1574_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1574_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1574_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_completed_
      -- 
    cpelement_group_1827 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1826);
      predecessors(1) <= cp_elements(1832);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1827)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1827),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1828 transition  bypass 
    -- predecessors 367 
    -- successors 1825 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1571_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1571_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1571_completed_
      -- 
    cp_elements(1828) <= cp_elements(367);
    -- CP-element group 1829 transition  output  bypass 
    -- predecessors 1825 
    -- successors 1830 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Sample/rr
      -- 
    cp_elements(1829) <= cp_elements(1825);
    rr_7651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1829), ack => binary_1573_inst_req_0); -- 
    -- CP-element group 1830 transition  input  no-bypass 
    -- predecessors 1829 
    -- successors 1826 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Sample/ra
      -- 
    ra_7652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1573_inst_ack_0, ack => cp_elements(1830)); -- 
    -- CP-element group 1831 transition  output  bypass 
    -- predecessors 1826 
    -- successors 1832 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Update/cr
      -- 
    cp_elements(1831) <= cp_elements(1826);
    cr_7656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1831), ack => binary_1573_inst_req_1); -- 
    -- CP-element group 1832 transition  input  no-bypass 
    -- predecessors 1831 
    -- successors 1827 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1573_complete_Update/ca
      -- 
    ca_7657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1573_inst_ack_1, ack => cp_elements(1832)); -- 
    -- CP-element group 1833 join  fork  transition  no-bypass 
    -- predecessors 1836 1837 
    -- successors 1834 1838 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_trigger_
      -- 
    cpelement_group_1833 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1836);
      predecessors(1) <= cp_elements(1837);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1833)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1833),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1834 join  fork  transition  no-bypass 
    -- predecessors 1833 1839 
    -- successors 1835 1840 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_active_
      -- 
    cpelement_group_1834 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1833);
      predecessors(1) <= cp_elements(1839);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1834)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1834),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1835 join  transition  bypass 
    -- predecessors 1834 1841 
    -- successors 1851 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1579_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1579_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1579_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1586_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1586_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1586_completed_
      -- 
    cpelement_group_1835 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1834);
      predecessors(1) <= cp_elements(1841);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1835)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1835),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1836 transition  bypass 
    -- predecessors 1729 
    -- successors 1833 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1576_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1576_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1576_completed_
      -- 
    cp_elements(1836) <= cp_elements(1729);
    -- CP-element group 1837 transition  bypass 
    -- predecessors 1114 
    -- successors 1833 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1577_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1577_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1577_completed_
      -- 
    cp_elements(1837) <= cp_elements(1114);
    -- CP-element group 1838 transition  output  bypass 
    -- predecessors 1833 
    -- successors 1839 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Sample/rr
      -- 
    cp_elements(1838) <= cp_elements(1833);
    rr_7673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1838), ack => binary_1578_inst_req_0); -- 
    -- CP-element group 1839 transition  input  no-bypass 
    -- predecessors 1838 
    -- successors 1834 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Sample/ra
      -- 
    ra_7674_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1578_inst_ack_0, ack => cp_elements(1839)); -- 
    -- CP-element group 1840 transition  output  bypass 
    -- predecessors 1834 
    -- successors 1841 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Update/cr
      -- 
    cp_elements(1840) <= cp_elements(1834);
    cr_7678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1840), ack => binary_1578_inst_req_1); -- 
    -- CP-element group 1841 transition  input  no-bypass 
    -- predecessors 1840 
    -- successors 1835 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1578_complete_Update/ca
      -- 
    ca_7679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1578_inst_ack_1, ack => cp_elements(1841)); -- 
    -- CP-element group 1842 join  fork  transition  no-bypass 
    -- predecessors 1845 1846 
    -- successors 1843 1847 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_trigger_
      -- 
    cpelement_group_1842 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1845);
      predecessors(1) <= cp_elements(1846);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1842)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1842),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1843 join  fork  transition  no-bypass 
    -- predecessors 1842 1848 
    -- successors 1844 1849 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_active_
      -- 
    cpelement_group_1843 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1842);
      predecessors(1) <= cp_elements(1848);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1843)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1843),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1844 join  transition  bypass 
    -- predecessors 1843 1850 
    -- successors 1851 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1584_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1584_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1584_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1587_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1587_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1587_completed_
      -- 
    cpelement_group_1844 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1843);
      predecessors(1) <= cp_elements(1850);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1844)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1844),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1845 transition  bypass 
    -- predecessors 1739 
    -- successors 1842 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1581_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1581_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1581_completed_
      -- 
    cp_elements(1845) <= cp_elements(1739);
    -- CP-element group 1846 transition  bypass 
    -- predecessors 1124 
    -- successors 1842 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1582_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1582_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1582_completed_
      -- 
    cp_elements(1846) <= cp_elements(1124);
    -- CP-element group 1847 transition  output  bypass 
    -- predecessors 1842 
    -- successors 1848 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Sample/rr
      -- 
    cp_elements(1847) <= cp_elements(1842);
    rr_7695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1847), ack => binary_1583_inst_req_0); -- 
    -- CP-element group 1848 transition  input  no-bypass 
    -- predecessors 1847 
    -- successors 1843 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Sample/ra
      -- 
    ra_7696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1583_inst_ack_0, ack => cp_elements(1848)); -- 
    -- CP-element group 1849 transition  output  bypass 
    -- predecessors 1843 
    -- successors 1850 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Update/cr
      -- 
    cp_elements(1849) <= cp_elements(1843);
    cr_7700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1849), ack => binary_1583_inst_req_1); -- 
    -- CP-element group 1850 transition  input  no-bypass 
    -- predecessors 1849 
    -- successors 1844 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1583_complete_Update/ca
      -- 
    ca_7701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1583_inst_ack_1, ack => cp_elements(1850)); -- 
    -- CP-element group 1851 join  fork  transition  bypass 
    -- predecessors 1835 1844 
    -- successors 1852 1854 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_trigger_
      -- 
    cpelement_group_1851 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1835);
      predecessors(1) <= cp_elements(1844);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1851)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1851),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1852 join  fork  transition  no-bypass 
    -- predecessors 1851 1855 
    -- successors 1853 1856 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_active_
      -- 
    cpelement_group_1852 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1851);
      predecessors(1) <= cp_elements(1855);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1852)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1852),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1853 join  transition  no-bypass 
    -- predecessors 1852 1857 
    -- successors 1883 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1589_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1589_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1589_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1606_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1606_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1606_completed_
      -- 
    cpelement_group_1853 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1852);
      predecessors(1) <= cp_elements(1857);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1853)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1853),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1854 transition  output  bypass 
    -- predecessors 1851 
    -- successors 1855 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Sample/rr
      -- 
    cp_elements(1854) <= cp_elements(1851);
    rr_7717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1854), ack => binary_1588_inst_req_0); -- 
    -- CP-element group 1855 transition  input  no-bypass 
    -- predecessors 1854 
    -- successors 1852 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Sample/ra
      -- 
    ra_7718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1588_inst_ack_0, ack => cp_elements(1855)); -- 
    -- CP-element group 1856 transition  output  bypass 
    -- predecessors 1852 
    -- successors 1857 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Update/cr
      -- 
    cp_elements(1856) <= cp_elements(1852);
    cr_7722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1856), ack => binary_1588_inst_req_1); -- 
    -- CP-element group 1857 transition  input  no-bypass 
    -- predecessors 1856 
    -- successors 1853 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1588_complete_Update/ca
      -- 
    ca_7723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1588_inst_ack_1, ack => cp_elements(1857)); -- 
    -- CP-element group 1858 join  fork  transition  no-bypass 
    -- predecessors 1861 1862 
    -- successors 1859 1863 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_trigger_
      -- 
    cpelement_group_1858 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1861);
      predecessors(1) <= cp_elements(1862);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1858)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1858),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1859 join  fork  transition  no-bypass 
    -- predecessors 1858 1864 
    -- successors 1860 1865 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_active_
      -- 
    cpelement_group_1859 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1858);
      predecessors(1) <= cp_elements(1864);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1859)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1859),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1860 join  transition  bypass 
    -- predecessors 1859 1866 
    -- successors 1876 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1594_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1594_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1594_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1601_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1601_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1601_completed_
      -- 
    cpelement_group_1860 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1859);
      predecessors(1) <= cp_elements(1866);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1860)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1860),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1861 transition  bypass 
    -- predecessors 1749 
    -- successors 1858 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1591_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1591_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1591_completed_
      -- 
    cp_elements(1861) <= cp_elements(1749);
    -- CP-element group 1862 transition  bypass 
    -- predecessors 1134 
    -- successors 1858 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1592_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1592_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1592_completed_
      -- 
    cp_elements(1862) <= cp_elements(1134);
    -- CP-element group 1863 transition  output  bypass 
    -- predecessors 1858 
    -- successors 1864 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Sample/rr
      -- 
    cp_elements(1863) <= cp_elements(1858);
    rr_7739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1863), ack => binary_1593_inst_req_0); -- 
    -- CP-element group 1864 transition  input  no-bypass 
    -- predecessors 1863 
    -- successors 1859 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Sample/ra
      -- 
    ra_7740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1593_inst_ack_0, ack => cp_elements(1864)); -- 
    -- CP-element group 1865 transition  output  bypass 
    -- predecessors 1859 
    -- successors 1866 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Update/cr
      -- 
    cp_elements(1865) <= cp_elements(1859);
    cr_7744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1865), ack => binary_1593_inst_req_1); -- 
    -- CP-element group 1866 transition  input  no-bypass 
    -- predecessors 1865 
    -- successors 1860 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1593_complete_Update/ca
      -- 
    ca_7745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1593_inst_ack_1, ack => cp_elements(1866)); -- 
    -- CP-element group 1867 join  fork  transition  no-bypass 
    -- predecessors 1870 1871 
    -- successors 1868 1872 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_trigger_
      -- 
    cpelement_group_1867 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1870);
      predecessors(1) <= cp_elements(1871);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1867)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1867),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1868 join  fork  transition  no-bypass 
    -- predecessors 1867 1873 
    -- successors 1869 1874 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_active_
      -- 
    cpelement_group_1868 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1867);
      predecessors(1) <= cp_elements(1873);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1868)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1868),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1869 join  transition  bypass 
    -- predecessors 1868 1875 
    -- successors 1876 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1599_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1599_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1599_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1602_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1602_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1602_completed_
      -- 
    cpelement_group_1869 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1868);
      predecessors(1) <= cp_elements(1875);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1869)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1869),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1870 transition  bypass 
    -- predecessors 1759 
    -- successors 1867 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1596_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1596_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1596_completed_
      -- 
    cp_elements(1870) <= cp_elements(1759);
    -- CP-element group 1871 transition  bypass 
    -- predecessors 1144 
    -- successors 1867 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1597_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1597_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1597_completed_
      -- 
    cp_elements(1871) <= cp_elements(1144);
    -- CP-element group 1872 transition  output  bypass 
    -- predecessors 1867 
    -- successors 1873 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Sample/rr
      -- 
    cp_elements(1872) <= cp_elements(1867);
    rr_7761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1872), ack => binary_1598_inst_req_0); -- 
    -- CP-element group 1873 transition  input  no-bypass 
    -- predecessors 1872 
    -- successors 1868 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Sample/ra
      -- 
    ra_7762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1598_inst_ack_0, ack => cp_elements(1873)); -- 
    -- CP-element group 1874 transition  output  bypass 
    -- predecessors 1868 
    -- successors 1875 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Update/cr
      -- 
    cp_elements(1874) <= cp_elements(1868);
    cr_7766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1874), ack => binary_1598_inst_req_1); -- 
    -- CP-element group 1875 transition  input  no-bypass 
    -- predecessors 1874 
    -- successors 1869 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1598_complete_Update/ca
      -- 
    ca_7767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1598_inst_ack_1, ack => cp_elements(1875)); -- 
    -- CP-element group 1876 join  fork  transition  bypass 
    -- predecessors 1860 1869 
    -- successors 1877 1879 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_trigger_
      -- 
    cpelement_group_1876 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1860);
      predecessors(1) <= cp_elements(1869);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1876)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1876),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1877 join  fork  transition  no-bypass 
    -- predecessors 1876 1880 
    -- successors 1878 1881 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_active_
      -- 
    cpelement_group_1877 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1876);
      predecessors(1) <= cp_elements(1880);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1877)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1877),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1878 join  transition  no-bypass 
    -- predecessors 1877 1882 
    -- successors 1883 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1604_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1604_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1604_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1607_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1607_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1607_completed_
      -- 
    cpelement_group_1878 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1877);
      predecessors(1) <= cp_elements(1882);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1878)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1878),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1879 transition  output  bypass 
    -- predecessors 1876 
    -- successors 1880 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Sample/rr
      -- 
    cp_elements(1879) <= cp_elements(1876);
    rr_7783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1879), ack => binary_1603_inst_req_0); -- 
    -- CP-element group 1880 transition  input  no-bypass 
    -- predecessors 1879 
    -- successors 1877 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Sample/ra
      -- 
    ra_7784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1603_inst_ack_0, ack => cp_elements(1880)); -- 
    -- CP-element group 1881 transition  output  bypass 
    -- predecessors 1877 
    -- successors 1882 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Update/cr
      -- 
    cp_elements(1881) <= cp_elements(1877);
    cr_7788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1881), ack => binary_1603_inst_req_1); -- 
    -- CP-element group 1882 transition  input  no-bypass 
    -- predecessors 1881 
    -- successors 1878 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1603_complete_Update/ca
      -- 
    ca_7789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1603_inst_ack_1, ack => cp_elements(1882)); -- 
    -- CP-element group 1883 join  fork  transition  bypass 
    -- predecessors 1853 1878 
    -- successors 1884 1886 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_trigger_
      -- 
    cpelement_group_1883 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1853);
      predecessors(1) <= cp_elements(1878);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1883)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1883),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1884 join  fork  transition  no-bypass 
    -- predecessors 1883 1887 
    -- successors 1885 1888 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_active_
      -- 
    cpelement_group_1884 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1883);
      predecessors(1) <= cp_elements(1887);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1884)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1884),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1885 join  transition  no-bypass 
    -- predecessors 1884 1889 
    -- successors 1890 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1609_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1609_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1609_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1612_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1612_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1612_completed_
      -- 
    cpelement_group_1885 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1884);
      predecessors(1) <= cp_elements(1889);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1885)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1885),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1886 transition  output  bypass 
    -- predecessors 1883 
    -- successors 1887 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Sample/rr
      -- 
    cp_elements(1886) <= cp_elements(1883);
    rr_7805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1886), ack => binary_1608_inst_req_0); -- 
    -- CP-element group 1887 transition  input  no-bypass 
    -- predecessors 1886 
    -- successors 1884 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Sample/ra
      -- 
    ra_7806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1608_inst_ack_0, ack => cp_elements(1887)); -- 
    -- CP-element group 1888 transition  output  bypass 
    -- predecessors 1884 
    -- successors 1889 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Update/cr
      -- 
    cp_elements(1888) <= cp_elements(1884);
    cr_7810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1888), ack => binary_1608_inst_req_1); -- 
    -- CP-element group 1889 transition  input  no-bypass 
    -- predecessors 1888 
    -- successors 1885 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1608_complete_Update/ca
      -- 
    ca_7811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1608_inst_ack_1, ack => cp_elements(1889)); -- 
    -- CP-element group 1890 join  fork  transition  no-bypass 
    -- predecessors 1885 1893 
    -- successors 1891 1894 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_trigger_
      -- 
    cpelement_group_1890 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1885);
      predecessors(1) <= cp_elements(1893);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1890)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1890),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1891 join  fork  transition  bypass 
    -- predecessors 1890 1895 
    -- successors 1892 1896 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_active_
      -- 
    cpelement_group_1891 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1890);
      predecessors(1) <= cp_elements(1895);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1891)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1891),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1892 join  transition  bypass 
    -- predecessors 1891 1897 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1614_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1614_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1614_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_completed_
      -- 
    cpelement_group_1892 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1891);
      predecessors(1) <= cp_elements(1897);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1892)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1892),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1893 transition  bypass 
    -- predecessors 367 
    -- successors 1890 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1611_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1611_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1611_completed_
      -- 
    cp_elements(1893) <= cp_elements(367);
    -- CP-element group 1894 transition  output  bypass 
    -- predecessors 1890 
    -- successors 1895 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Sample/rr
      -- 
    cp_elements(1894) <= cp_elements(1890);
    rr_7827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1894), ack => binary_1613_inst_req_0); -- 
    -- CP-element group 1895 transition  input  no-bypass 
    -- predecessors 1894 
    -- successors 1891 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Sample/ra
      -- 
    ra_7828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1613_inst_ack_0, ack => cp_elements(1895)); -- 
    -- CP-element group 1896 transition  output  bypass 
    -- predecessors 1891 
    -- successors 1897 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Update/cr
      -- 
    cp_elements(1896) <= cp_elements(1891);
    cr_7832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1896), ack => binary_1613_inst_req_1); -- 
    -- CP-element group 1897 transition  input  no-bypass 
    -- predecessors 1896 
    -- successors 1892 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1613_complete_Update/ca
      -- 
    ca_7833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1613_inst_ack_1, ack => cp_elements(1897)); -- 
    -- CP-element group 1898 join  fork  transition  no-bypass 
    -- predecessors 1901 1902 
    -- successors 1899 1903 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_trigger_
      -- 
    cpelement_group_1898 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1901);
      predecessors(1) <= cp_elements(1902);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1898)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1898),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1899 join  fork  transition  no-bypass 
    -- predecessors 1898 1904 
    -- successors 1900 1905 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_active_
      -- 
    cpelement_group_1899 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1898);
      predecessors(1) <= cp_elements(1904);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1899)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1899),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1900 join  transition  bypass 
    -- predecessors 1899 1906 
    -- successors 1916 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1619_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1619_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1619_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1626_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1626_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1626_completed_
      -- 
    cpelement_group_1900 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1899);
      predecessors(1) <= cp_elements(1906);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1900)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1900),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1901 transition  bypass 
    -- predecessors 1729 
    -- successors 1898 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1616_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1616_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1616_completed_
      -- 
    cp_elements(1901) <= cp_elements(1729);
    -- CP-element group 1902 transition  bypass 
    -- predecessors 1219 
    -- successors 1898 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1617_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1617_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1617_completed_
      -- 
    cp_elements(1902) <= cp_elements(1219);
    -- CP-element group 1903 transition  output  bypass 
    -- predecessors 1898 
    -- successors 1904 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Sample/rr
      -- 
    cp_elements(1903) <= cp_elements(1898);
    rr_7849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1903), ack => binary_1618_inst_req_0); -- 
    -- CP-element group 1904 transition  input  no-bypass 
    -- predecessors 1903 
    -- successors 1899 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Sample/ra
      -- 
    ra_7850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1618_inst_ack_0, ack => cp_elements(1904)); -- 
    -- CP-element group 1905 transition  output  bypass 
    -- predecessors 1899 
    -- successors 1906 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Update/cr
      -- 
    cp_elements(1905) <= cp_elements(1899);
    cr_7854_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1905), ack => binary_1618_inst_req_1); -- 
    -- CP-element group 1906 transition  input  no-bypass 
    -- predecessors 1905 
    -- successors 1900 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1618_complete_Update/ca
      -- 
    ca_7855_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1618_inst_ack_1, ack => cp_elements(1906)); -- 
    -- CP-element group 1907 join  fork  transition  no-bypass 
    -- predecessors 1910 1911 
    -- successors 1908 1912 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_trigger_
      -- 
    cpelement_group_1907 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1910);
      predecessors(1) <= cp_elements(1911);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1907)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1907),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1908 join  fork  transition  no-bypass 
    -- predecessors 1907 1913 
    -- successors 1909 1914 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_active_
      -- 
    cpelement_group_1908 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1907);
      predecessors(1) <= cp_elements(1913);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1908)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1908),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1909 join  transition  bypass 
    -- predecessors 1908 1915 
    -- successors 1916 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1624_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1624_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1624_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1627_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1627_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1627_completed_
      -- 
    cpelement_group_1909 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1908);
      predecessors(1) <= cp_elements(1915);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1909)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1909),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1910 transition  bypass 
    -- predecessors 1739 
    -- successors 1907 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1621_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1621_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1621_completed_
      -- 
    cp_elements(1910) <= cp_elements(1739);
    -- CP-element group 1911 transition  bypass 
    -- predecessors 1229 
    -- successors 1907 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1622_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1622_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1622_completed_
      -- 
    cp_elements(1911) <= cp_elements(1229);
    -- CP-element group 1912 transition  output  bypass 
    -- predecessors 1907 
    -- successors 1913 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Sample/rr
      -- 
    cp_elements(1912) <= cp_elements(1907);
    rr_7871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1912), ack => binary_1623_inst_req_0); -- 
    -- CP-element group 1913 transition  input  no-bypass 
    -- predecessors 1912 
    -- successors 1908 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Sample/ra
      -- 
    ra_7872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1623_inst_ack_0, ack => cp_elements(1913)); -- 
    -- CP-element group 1914 transition  output  bypass 
    -- predecessors 1908 
    -- successors 1915 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Update/cr
      -- 
    cp_elements(1914) <= cp_elements(1908);
    cr_7876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1914), ack => binary_1623_inst_req_1); -- 
    -- CP-element group 1915 transition  input  no-bypass 
    -- predecessors 1914 
    -- successors 1909 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1623_complete_Update/ca
      -- 
    ca_7877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1623_inst_ack_1, ack => cp_elements(1915)); -- 
    -- CP-element group 1916 join  fork  transition  bypass 
    -- predecessors 1900 1909 
    -- successors 1917 1919 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_trigger_
      -- 
    cpelement_group_1916 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1900);
      predecessors(1) <= cp_elements(1909);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1916)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1916),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1917 join  fork  transition  no-bypass 
    -- predecessors 1916 1920 
    -- successors 1918 1921 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_active_
      -- 
    cpelement_group_1917 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1916);
      predecessors(1) <= cp_elements(1920);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1917)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1917),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1918 join  transition  no-bypass 
    -- predecessors 1917 1922 
    -- successors 1948 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1646_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1646_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1646_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1629_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1629_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1629_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_completed_
      -- 
    cpelement_group_1918 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1917);
      predecessors(1) <= cp_elements(1922);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1918)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1918),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1919 transition  output  bypass 
    -- predecessors 1916 
    -- successors 1920 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Sample/rr
      -- 
    cp_elements(1919) <= cp_elements(1916);
    rr_7893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1919), ack => binary_1628_inst_req_0); -- 
    -- CP-element group 1920 transition  input  no-bypass 
    -- predecessors 1919 
    -- successors 1917 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Sample/ra
      -- 
    ra_7894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1628_inst_ack_0, ack => cp_elements(1920)); -- 
    -- CP-element group 1921 transition  output  bypass 
    -- predecessors 1917 
    -- successors 1922 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Update/cr
      -- 
    cp_elements(1921) <= cp_elements(1917);
    cr_7898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1921), ack => binary_1628_inst_req_1); -- 
    -- CP-element group 1922 transition  input  no-bypass 
    -- predecessors 1921 
    -- successors 1918 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1628_complete_Update/ca
      -- 
    ca_7899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1628_inst_ack_1, ack => cp_elements(1922)); -- 
    -- CP-element group 1923 join  fork  transition  no-bypass 
    -- predecessors 1926 1927 
    -- successors 1924 1928 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_trigger_
      -- 
    cpelement_group_1923 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1926);
      predecessors(1) <= cp_elements(1927);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1923)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1923),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1924 join  fork  transition  no-bypass 
    -- predecessors 1923 1929 
    -- successors 1925 1930 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_active_
      -- 
    cpelement_group_1924 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1923);
      predecessors(1) <= cp_elements(1929);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1924)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1924),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1925 join  transition  bypass 
    -- predecessors 1924 1931 
    -- successors 1941 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1641_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1641_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1641_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1634_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1634_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1634_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_completed_
      -- 
    cpelement_group_1925 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1924);
      predecessors(1) <= cp_elements(1931);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1925)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1925),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1926 transition  bypass 
    -- predecessors 1749 
    -- successors 1923 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1631_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1631_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1631_completed_
      -- 
    cp_elements(1926) <= cp_elements(1749);
    -- CP-element group 1927 transition  bypass 
    -- predecessors 1239 
    -- successors 1923 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1632_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1632_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1632_completed_
      -- 
    cp_elements(1927) <= cp_elements(1239);
    -- CP-element group 1928 transition  output  bypass 
    -- predecessors 1923 
    -- successors 1929 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Sample/rr
      -- 
    cp_elements(1928) <= cp_elements(1923);
    rr_7915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1928), ack => binary_1633_inst_req_0); -- 
    -- CP-element group 1929 transition  input  no-bypass 
    -- predecessors 1928 
    -- successors 1924 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Sample/ra
      -- 
    ra_7916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1633_inst_ack_0, ack => cp_elements(1929)); -- 
    -- CP-element group 1930 transition  output  bypass 
    -- predecessors 1924 
    -- successors 1931 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Update/$entry
      -- 
    cp_elements(1930) <= cp_elements(1924);
    cr_7920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1930), ack => binary_1633_inst_req_1); -- 
    -- CP-element group 1931 transition  input  no-bypass 
    -- predecessors 1930 
    -- successors 1925 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1633_complete_Update/ca
      -- 
    ca_7921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1633_inst_ack_1, ack => cp_elements(1931)); -- 
    -- CP-element group 1932 join  fork  transition  no-bypass 
    -- predecessors 1935 1936 
    -- successors 1933 1937 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_trigger_
      -- 
    cpelement_group_1932 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1935);
      predecessors(1) <= cp_elements(1936);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1932)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1932),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1933 join  fork  transition  no-bypass 
    -- predecessors 1932 1938 
    -- successors 1934 1939 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_active_
      -- 
    cpelement_group_1933 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1932);
      predecessors(1) <= cp_elements(1938);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1933)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1933),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1934 join  transition  bypass 
    -- predecessors 1933 1940 
    -- successors 1941 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1639_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1639_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1639_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1642_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1642_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1642_completed_
      -- 
    cpelement_group_1934 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1933);
      predecessors(1) <= cp_elements(1940);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1934)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1934),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1935 transition  bypass 
    -- predecessors 1759 
    -- successors 1932 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1636_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1636_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1636_completed_
      -- 
    cp_elements(1935) <= cp_elements(1759);
    -- CP-element group 1936 transition  bypass 
    -- predecessors 1249 
    -- successors 1932 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1637_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1637_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1637_completed_
      -- 
    cp_elements(1936) <= cp_elements(1249);
    -- CP-element group 1937 transition  output  bypass 
    -- predecessors 1932 
    -- successors 1938 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Sample/rr
      -- 
    cp_elements(1937) <= cp_elements(1932);
    rr_7937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1937), ack => binary_1638_inst_req_0); -- 
    -- CP-element group 1938 transition  input  no-bypass 
    -- predecessors 1937 
    -- successors 1933 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Sample/ra
      -- 
    ra_7938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1638_inst_ack_0, ack => cp_elements(1938)); -- 
    -- CP-element group 1939 transition  output  bypass 
    -- predecessors 1933 
    -- successors 1940 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Update/cr
      -- 
    cp_elements(1939) <= cp_elements(1933);
    cr_7942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1939), ack => binary_1638_inst_req_1); -- 
    -- CP-element group 1940 transition  input  no-bypass 
    -- predecessors 1939 
    -- successors 1934 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1638_complete_Update/ca
      -- 
    ca_7943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1638_inst_ack_1, ack => cp_elements(1940)); -- 
    -- CP-element group 1941 join  fork  transition  bypass 
    -- predecessors 1925 1934 
    -- successors 1942 1944 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_trigger_
      -- 
    cpelement_group_1941 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1925);
      predecessors(1) <= cp_elements(1934);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1941)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1941),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1942 join  fork  transition  no-bypass 
    -- predecessors 1941 1945 
    -- successors 1943 1946 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_active_
      -- 
    cpelement_group_1942 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1941);
      predecessors(1) <= cp_elements(1945);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1942)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1942),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1943 join  transition  no-bypass 
    -- predecessors 1942 1947 
    -- successors 1948 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1644_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1647_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1644_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1644_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1647_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1647_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_completed_
      -- 
    cpelement_group_1943 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1942);
      predecessors(1) <= cp_elements(1947);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1943)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1943),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1944 transition  output  bypass 
    -- predecessors 1941 
    -- successors 1945 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Sample/$entry
      -- 
    cp_elements(1944) <= cp_elements(1941);
    rr_7959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1944), ack => binary_1643_inst_req_0); -- 
    -- CP-element group 1945 transition  input  no-bypass 
    -- predecessors 1944 
    -- successors 1942 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Sample/ra
      -- 
    ra_7960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1643_inst_ack_0, ack => cp_elements(1945)); -- 
    -- CP-element group 1946 transition  output  bypass 
    -- predecessors 1942 
    -- successors 1947 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Update/cr
      -- 
    cp_elements(1946) <= cp_elements(1942);
    cr_7964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1946), ack => binary_1643_inst_req_1); -- 
    -- CP-element group 1947 transition  input  no-bypass 
    -- predecessors 1946 
    -- successors 1943 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1643_complete_Update/ca
      -- 
    ca_7965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1643_inst_ack_1, ack => cp_elements(1947)); -- 
    -- CP-element group 1948 join  fork  transition  bypass 
    -- predecessors 1918 1943 
    -- successors 1949 1951 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_trigger_
      -- 
    cpelement_group_1948 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1918);
      predecessors(1) <= cp_elements(1943);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1948)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1948),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1949 join  fork  transition  no-bypass 
    -- predecessors 1948 1952 
    -- successors 1950 1953 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_active_
      -- 
    cpelement_group_1949 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1948);
      predecessors(1) <= cp_elements(1952);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1949)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1949),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1950 join  transition  no-bypass 
    -- predecessors 1949 1954 
    -- successors 1955 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1649_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1649_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1649_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1652_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1652_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1652_completed_
      -- 
    cpelement_group_1950 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1949);
      predecessors(1) <= cp_elements(1954);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1950)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1950),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1951 transition  output  bypass 
    -- predecessors 1948 
    -- successors 1952 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Sample/rr
      -- 
    cp_elements(1951) <= cp_elements(1948);
    rr_7981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1951), ack => binary_1648_inst_req_0); -- 
    -- CP-element group 1952 transition  input  no-bypass 
    -- predecessors 1951 
    -- successors 1949 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Sample/ra
      -- 
    ra_7982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1648_inst_ack_0, ack => cp_elements(1952)); -- 
    -- CP-element group 1953 transition  output  bypass 
    -- predecessors 1949 
    -- successors 1954 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Update/cr
      -- 
    cp_elements(1953) <= cp_elements(1949);
    cr_7986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1953), ack => binary_1648_inst_req_1); -- 
    -- CP-element group 1954 transition  input  no-bypass 
    -- predecessors 1953 
    -- successors 1950 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1648_complete_Update/ca
      -- 
    ca_7987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1648_inst_ack_1, ack => cp_elements(1954)); -- 
    -- CP-element group 1955 join  fork  transition  no-bypass 
    -- predecessors 1950 1958 
    -- successors 1956 1959 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_trigger_
      -- 
    cpelement_group_1955 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1950);
      predecessors(1) <= cp_elements(1958);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1955)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1955),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1956 join  fork  transition  bypass 
    -- predecessors 1955 1960 
    -- successors 1957 1961 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_active_
      -- 
    cpelement_group_1956 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1955);
      predecessors(1) <= cp_elements(1960);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1956)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1956),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1957 join  transition  bypass 
    -- predecessors 1956 1962 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1654_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1654_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1654_completed_
      -- 
    cpelement_group_1957 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1956);
      predecessors(1) <= cp_elements(1962);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1957)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1957),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1958 transition  bypass 
    -- predecessors 367 
    -- successors 1955 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1651_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1651_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1651_completed_
      -- 
    cp_elements(1958) <= cp_elements(367);
    -- CP-element group 1959 transition  output  bypass 
    -- predecessors 1955 
    -- successors 1960 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Sample/rr
      -- 
    cp_elements(1959) <= cp_elements(1955);
    rr_8003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1959), ack => binary_1653_inst_req_0); -- 
    -- CP-element group 1960 transition  input  no-bypass 
    -- predecessors 1959 
    -- successors 1956 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Sample/ra
      -- 
    ra_8004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1653_inst_ack_0, ack => cp_elements(1960)); -- 
    -- CP-element group 1961 transition  output  bypass 
    -- predecessors 1956 
    -- successors 1962 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Update/$entry
      -- 
    cp_elements(1961) <= cp_elements(1956);
    cr_8008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1961), ack => binary_1653_inst_req_1); -- 
    -- CP-element group 1962 transition  input  no-bypass 
    -- predecessors 1961 
    -- successors 1957 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1653_complete_Update/$exit
      -- 
    ca_8009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1653_inst_ack_1, ack => cp_elements(1962)); -- 
    -- CP-element group 1963 join  fork  transition  no-bypass 
    -- predecessors 1966 1967 
    -- successors 1964 1968 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_trigger_
      -- 
    cpelement_group_1963 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1966);
      predecessors(1) <= cp_elements(1967);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1963)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1963),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1964 join  fork  transition  no-bypass 
    -- predecessors 1963 1969 
    -- successors 1965 1970 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_active_
      -- 
    cpelement_group_1964 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1963);
      predecessors(1) <= cp_elements(1969);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1964)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1964),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1965 join  transition  bypass 
    -- predecessors 1964 1971 
    -- successors 1981 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1659_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1659_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1666_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1666_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1659_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1666_trigger_
      -- 
    cpelement_group_1965 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1964);
      predecessors(1) <= cp_elements(1971);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1965)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1965),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1966 transition  bypass 
    -- predecessors 1729 
    -- successors 1963 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1656_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1656_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1656_trigger_
      -- 
    cp_elements(1966) <= cp_elements(1729);
    -- CP-element group 1967 transition  bypass 
    -- predecessors 1324 
    -- successors 1963 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1657_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1657_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1657_completed_
      -- 
    cp_elements(1967) <= cp_elements(1324);
    -- CP-element group 1968 transition  output  bypass 
    -- predecessors 1963 
    -- successors 1969 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Sample/$entry
      -- 
    cp_elements(1968) <= cp_elements(1963);
    rr_8025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1968), ack => binary_1658_inst_req_0); -- 
    -- CP-element group 1969 transition  input  no-bypass 
    -- predecessors 1968 
    -- successors 1964 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Sample/$exit
      -- 
    ra_8026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1658_inst_ack_0, ack => cp_elements(1969)); -- 
    -- CP-element group 1970 transition  output  bypass 
    -- predecessors 1964 
    -- successors 1971 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Update/$entry
      -- 
    cp_elements(1970) <= cp_elements(1964);
    cr_8030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1970), ack => binary_1658_inst_req_1); -- 
    -- CP-element group 1971 transition  input  no-bypass 
    -- predecessors 1970 
    -- successors 1965 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1658_complete_Update/ca
      -- 
    ca_8031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1658_inst_ack_1, ack => cp_elements(1971)); -- 
    -- CP-element group 1972 join  fork  transition  no-bypass 
    -- predecessors 1975 1976 
    -- successors 1973 1977 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_trigger_
      -- 
    cpelement_group_1972 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1975);
      predecessors(1) <= cp_elements(1976);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1972)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1972),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1973 join  fork  transition  no-bypass 
    -- predecessors 1972 1978 
    -- successors 1974 1979 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_active_
      -- 
    cpelement_group_1973 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1972);
      predecessors(1) <= cp_elements(1978);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1973)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1973),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1974 join  transition  bypass 
    -- predecessors 1973 1980 
    -- successors 1981 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1667_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1667_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1667_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1664_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1664_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1664_completed_
      -- 
    cpelement_group_1974 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1973);
      predecessors(1) <= cp_elements(1980);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1974)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1974),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1975 transition  bypass 
    -- predecessors 1739 
    -- successors 1972 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1661_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1661_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1661_trigger_
      -- 
    cp_elements(1975) <= cp_elements(1739);
    -- CP-element group 1976 transition  bypass 
    -- predecessors 1334 
    -- successors 1972 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1662_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1662_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1662_completed_
      -- 
    cp_elements(1976) <= cp_elements(1334);
    -- CP-element group 1977 transition  output  bypass 
    -- predecessors 1972 
    -- successors 1978 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Sample/rr
      -- 
    cp_elements(1977) <= cp_elements(1972);
    rr_8047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1977), ack => binary_1663_inst_req_0); -- 
    -- CP-element group 1978 transition  input  no-bypass 
    -- predecessors 1977 
    -- successors 1973 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Sample/$exit
      -- 
    ra_8048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1663_inst_ack_0, ack => cp_elements(1978)); -- 
    -- CP-element group 1979 transition  output  bypass 
    -- predecessors 1973 
    -- successors 1980 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Update/cr
      -- 
    cp_elements(1979) <= cp_elements(1973);
    cr_8052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1979), ack => binary_1663_inst_req_1); -- 
    -- CP-element group 1980 transition  input  no-bypass 
    -- predecessors 1979 
    -- successors 1974 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1663_complete_Update/ca
      -- 
    ca_8053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1663_inst_ack_1, ack => cp_elements(1980)); -- 
    -- CP-element group 1981 join  fork  transition  bypass 
    -- predecessors 1965 1974 
    -- successors 1982 1984 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_trigger_
      -- 
    cpelement_group_1981 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1965);
      predecessors(1) <= cp_elements(1974);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1981)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1981),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1982 join  fork  transition  no-bypass 
    -- predecessors 1981 1985 
    -- successors 1983 1986 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_active_
      -- 
    cpelement_group_1982 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1981);
      predecessors(1) <= cp_elements(1985);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1982)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1982),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1983 join  transition  no-bypass 
    -- predecessors 1982 1987 
    -- successors 2013 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1669_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1669_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1669_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1686_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1686_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1686_completed_
      -- 
    cpelement_group_1983 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1982);
      predecessors(1) <= cp_elements(1987);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1983)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1983),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1984 transition  output  bypass 
    -- predecessors 1981 
    -- successors 1985 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Sample/rr
      -- 
    cp_elements(1984) <= cp_elements(1981);
    rr_8069_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1984), ack => binary_1668_inst_req_0); -- 
    -- CP-element group 1985 transition  input  no-bypass 
    -- predecessors 1984 
    -- successors 1982 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Sample/ra
      -- 
    ra_8070_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1668_inst_ack_0, ack => cp_elements(1985)); -- 
    -- CP-element group 1986 transition  output  bypass 
    -- predecessors 1982 
    -- successors 1987 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Update/cr
      -- 
    cp_elements(1986) <= cp_elements(1982);
    cr_8074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1986), ack => binary_1668_inst_req_1); -- 
    -- CP-element group 1987 transition  input  no-bypass 
    -- predecessors 1986 
    -- successors 1983 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1668_complete_Update/ca
      -- 
    ca_8075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1668_inst_ack_1, ack => cp_elements(1987)); -- 
    -- CP-element group 1988 join  fork  transition  no-bypass 
    -- predecessors 1991 1992 
    -- successors 1989 1993 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_trigger_
      -- 
    cpelement_group_1988 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1991);
      predecessors(1) <= cp_elements(1992);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1988)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1988),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1989 join  fork  transition  no-bypass 
    -- predecessors 1988 1994 
    -- successors 1990 1995 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_active_
      -- 
    cpelement_group_1989 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1988);
      predecessors(1) <= cp_elements(1994);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1989)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1989),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1990 join  transition  bypass 
    -- predecessors 1989 1996 
    -- successors 2006 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1674_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1674_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1674_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1681_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1681_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1681_completed_
      -- 
    cpelement_group_1990 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1989);
      predecessors(1) <= cp_elements(1996);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1990)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1990),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1991 transition  bypass 
    -- predecessors 1749 
    -- successors 1988 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1671_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1671_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1671_completed_
      -- 
    cp_elements(1991) <= cp_elements(1749);
    -- CP-element group 1992 transition  bypass 
    -- predecessors 1344 
    -- successors 1988 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1672_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1672_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1672_completed_
      -- 
    cp_elements(1992) <= cp_elements(1344);
    -- CP-element group 1993 transition  output  bypass 
    -- predecessors 1988 
    -- successors 1994 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Sample/rr
      -- 
    cp_elements(1993) <= cp_elements(1988);
    rr_8091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1993), ack => binary_1673_inst_req_0); -- 
    -- CP-element group 1994 transition  input  no-bypass 
    -- predecessors 1993 
    -- successors 1989 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Sample/ra
      -- 
    ra_8092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1673_inst_ack_0, ack => cp_elements(1994)); -- 
    -- CP-element group 1995 transition  output  bypass 
    -- predecessors 1989 
    -- successors 1996 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Update/cr
      -- 
    cp_elements(1995) <= cp_elements(1989);
    cr_8096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1995), ack => binary_1673_inst_req_1); -- 
    -- CP-element group 1996 transition  input  no-bypass 
    -- predecessors 1995 
    -- successors 1990 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1673_complete_Update/ca
      -- 
    ca_8097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1673_inst_ack_1, ack => cp_elements(1996)); -- 
    -- CP-element group 1997 join  fork  transition  no-bypass 
    -- predecessors 2000 2001 
    -- successors 1998 2002 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_trigger_
      -- 
    cpelement_group_1997 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2000);
      predecessors(1) <= cp_elements(2001);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1997)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1997),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1998 join  fork  transition  no-bypass 
    -- predecessors 1997 2003 
    -- successors 1999 2004 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_active_
      -- 
    cpelement_group_1998 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1997);
      predecessors(1) <= cp_elements(2003);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(1998)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1998),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1999 join  transition  bypass 
    -- predecessors 1998 2005 
    -- successors 2006 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1679_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1679_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1679_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1682_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1682_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1682_completed_
      -- 
    cpelement_group_1999 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1998);
      predecessors(1) <= cp_elements(2005);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(1999)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1999),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2000 transition  bypass 
    -- predecessors 1759 
    -- successors 1997 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1676_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1676_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1676_completed_
      -- 
    cp_elements(2000) <= cp_elements(1759);
    -- CP-element group 2001 transition  bypass 
    -- predecessors 1354 
    -- successors 1997 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1677_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1677_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1677_completed_
      -- 
    cp_elements(2001) <= cp_elements(1354);
    -- CP-element group 2002 transition  output  bypass 
    -- predecessors 1997 
    -- successors 2003 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Sample/rr
      -- 
    cp_elements(2002) <= cp_elements(1997);
    rr_8113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2002), ack => binary_1678_inst_req_0); -- 
    -- CP-element group 2003 transition  input  no-bypass 
    -- predecessors 2002 
    -- successors 1998 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Sample/ra
      -- 
    ra_8114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1678_inst_ack_0, ack => cp_elements(2003)); -- 
    -- CP-element group 2004 transition  output  bypass 
    -- predecessors 1998 
    -- successors 2005 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Update/cr
      -- 
    cp_elements(2004) <= cp_elements(1998);
    cr_8118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2004), ack => binary_1678_inst_req_1); -- 
    -- CP-element group 2005 transition  input  no-bypass 
    -- predecessors 2004 
    -- successors 1999 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1678_complete_Update/ca
      -- 
    ca_8119_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1678_inst_ack_1, ack => cp_elements(2005)); -- 
    -- CP-element group 2006 join  fork  transition  bypass 
    -- predecessors 1990 1999 
    -- successors 2007 2009 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_trigger_
      -- 
    cpelement_group_2006 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1990);
      predecessors(1) <= cp_elements(1999);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2006)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2006),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2007 join  fork  transition  no-bypass 
    -- predecessors 2006 2010 
    -- successors 2008 2011 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_active_
      -- 
    cpelement_group_2007 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2006);
      predecessors(1) <= cp_elements(2010);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2007)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2007),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2008 join  transition  no-bypass 
    -- predecessors 2007 2012 
    -- successors 2013 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1684_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1684_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1684_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1687_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1687_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1687_completed_
      -- 
    cpelement_group_2008 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2007);
      predecessors(1) <= cp_elements(2012);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2008)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2008),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2009 transition  output  bypass 
    -- predecessors 2006 
    -- successors 2010 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Sample/rr
      -- 
    cp_elements(2009) <= cp_elements(2006);
    rr_8135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2009), ack => binary_1683_inst_req_0); -- 
    -- CP-element group 2010 transition  input  no-bypass 
    -- predecessors 2009 
    -- successors 2007 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Sample/ra
      -- 
    ra_8136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1683_inst_ack_0, ack => cp_elements(2010)); -- 
    -- CP-element group 2011 transition  output  bypass 
    -- predecessors 2007 
    -- successors 2012 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Update/cr
      -- 
    cp_elements(2011) <= cp_elements(2007);
    cr_8140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2011), ack => binary_1683_inst_req_1); -- 
    -- CP-element group 2012 transition  input  no-bypass 
    -- predecessors 2011 
    -- successors 2008 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1683_complete_Update/ca
      -- 
    ca_8141_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1683_inst_ack_1, ack => cp_elements(2012)); -- 
    -- CP-element group 2013 join  fork  transition  bypass 
    -- predecessors 1983 2008 
    -- successors 2014 2016 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_trigger_
      -- 
    cpelement_group_2013 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1983);
      predecessors(1) <= cp_elements(2008);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2013)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2013),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2014 join  fork  transition  no-bypass 
    -- predecessors 2013 2017 
    -- successors 2015 2018 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_active_
      -- 
    cpelement_group_2014 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2013);
      predecessors(1) <= cp_elements(2017);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2014)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2014),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2015 join  transition  no-bypass 
    -- predecessors 2014 2019 
    -- successors 2020 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1689_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1689_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1689_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1692_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1692_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1692_completed_
      -- 
    cpelement_group_2015 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2014);
      predecessors(1) <= cp_elements(2019);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2015)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2015),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2016 transition  output  bypass 
    -- predecessors 2013 
    -- successors 2017 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Sample/rr
      -- 
    cp_elements(2016) <= cp_elements(2013);
    rr_8157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2016), ack => binary_1688_inst_req_0); -- 
    -- CP-element group 2017 transition  input  no-bypass 
    -- predecessors 2016 
    -- successors 2014 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Sample/ra
      -- 
    ra_8158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1688_inst_ack_0, ack => cp_elements(2017)); -- 
    -- CP-element group 2018 transition  output  bypass 
    -- predecessors 2014 
    -- successors 2019 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Update/cr
      -- 
    cp_elements(2018) <= cp_elements(2014);
    cr_8162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2018), ack => binary_1688_inst_req_1); -- 
    -- CP-element group 2019 transition  input  no-bypass 
    -- predecessors 2018 
    -- successors 2015 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1688_complete_Update/ca
      -- 
    ca_8163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1688_inst_ack_1, ack => cp_elements(2019)); -- 
    -- CP-element group 2020 join  fork  transition  no-bypass 
    -- predecessors 2015 2023 
    -- successors 2021 2024 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_trigger_
      -- 
    cpelement_group_2020 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2015);
      predecessors(1) <= cp_elements(2023);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2020)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2020),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2021 join  fork  transition  bypass 
    -- predecessors 2020 2025 
    -- successors 2022 2026 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_active_
      -- 
    cpelement_group_2021 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2020);
      predecessors(1) <= cp_elements(2025);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2021)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2021),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2022 join  transition  bypass 
    -- predecessors 2021 2027 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1694_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1694_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1694_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_completed_
      -- 
    cpelement_group_2022 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2021);
      predecessors(1) <= cp_elements(2027);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2022)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2022),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2023 transition  bypass 
    -- predecessors 367 
    -- successors 2020 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1691_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1691_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1691_completed_
      -- 
    cp_elements(2023) <= cp_elements(367);
    -- CP-element group 2024 transition  output  bypass 
    -- predecessors 2020 
    -- successors 2025 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Sample/rr
      -- 
    cp_elements(2024) <= cp_elements(2020);
    rr_8179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2024), ack => binary_1693_inst_req_0); -- 
    -- CP-element group 2025 transition  input  no-bypass 
    -- predecessors 2024 
    -- successors 2021 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Sample/ra
      -- 
    ra_8180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1693_inst_ack_0, ack => cp_elements(2025)); -- 
    -- CP-element group 2026 transition  output  bypass 
    -- predecessors 2021 
    -- successors 2027 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Update/cr
      -- 
    cp_elements(2026) <= cp_elements(2021);
    cr_8184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2026), ack => binary_1693_inst_req_1); -- 
    -- CP-element group 2027 transition  input  no-bypass 
    -- predecessors 2026 
    -- successors 2022 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1693_complete_Update/ca
      -- 
    ca_8185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1693_inst_ack_1, ack => cp_elements(2027)); -- 
    -- CP-element group 2028 join  fork  transition  bypass 
    -- predecessors 2032 2034 
    -- successors 2029 2035 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_active_
      -- 
    cpelement_group_2028 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2032);
      predecessors(1) <= cp_elements(2034);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2028)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2028),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2029 join  fork  transition  bypass 
    -- predecessors 2028 2037 
    -- successors 2071 2136 2201 2266 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1698_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1698_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1698_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_completed_
      -- 
    cpelement_group_2029 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2028);
      predecessors(1) <= cp_elements(2037);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2029)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2029),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2030 transition  input  output  no-bypass 
    -- predecessors 442 
    -- successors 2031 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8203_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1697_base_resize_ack_0, ack => cp_elements(2030)); -- 
    sum_rename_req_8207_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2030), ack => ptr_deref_1697_root_address_inst_req_0); -- 
    -- CP-element group 2031 transition  input  output  no-bypass 
    -- predecessors 2030 
    -- successors 2032 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8208_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1697_root_address_inst_ack_0, ack => cp_elements(2031)); -- 
    root_register_req_8212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2031), ack => ptr_deref_1697_addr_0_req_0); -- 
    -- CP-element group 2032 fork  transition  input  no-bypass 
    -- predecessors 2031 
    -- successors 2028 2033 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_word_addrgen/root_register_ack
      -- 
    root_register_ack_8213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1697_addr_0_ack_0, ack => cp_elements(2032)); -- 
    -- CP-element group 2033 transition  output  bypass 
    -- predecessors 2032 
    -- successors 2034 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/word_access/word_access_0/rr
      -- 
    cp_elements(2033) <= cp_elements(2032);
    rr_8223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2033), ack => ptr_deref_1697_load_0_req_0); -- 
    -- CP-element group 2034 transition  input  no-bypass 
    -- predecessors 2033 
    -- successors 2028 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_request/word_access/word_access_0/ra
      -- 
    ra_8224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1697_load_0_ack_0, ack => cp_elements(2034)); -- 
    -- CP-element group 2035 transition  output  bypass 
    -- predecessors 2028 
    -- successors 2036 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2035) <= cp_elements(2028);
    cr_8234_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2035), ack => ptr_deref_1697_load_0_req_1); -- 
    -- CP-element group 2036 transition  input  output  no-bypass 
    -- predecessors 2035 
    -- successors 2037 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/merge_req
      -- 
    ca_8235_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1697_load_0_ack_1, ack => cp_elements(2036)); -- 
    merge_req_8236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2036), ack => ptr_deref_1697_gather_scatter_req_0); -- 
    -- CP-element group 2037 transition  input  no-bypass 
    -- predecessors 2036 
    -- successors 2029 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1697_complete/merge_ack
      -- 
    merge_ack_8237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1697_gather_scatter_ack_0, ack => cp_elements(2037)); -- 
    -- CP-element group 2038 join  fork  transition  bypass 
    -- predecessors 2042 2044 
    -- successors 2039 2045 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_active_
      -- 
    cpelement_group_2038 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2042);
      predecessors(1) <= cp_elements(2044);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2038)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2038),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2039 join  fork  transition  bypass 
    -- predecessors 2038 2047 
    -- successors 2080 2145 2210 2275 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1702_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1702_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1702_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_completed_
      -- 
    cpelement_group_2039 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2038);
      predecessors(1) <= cp_elements(2047);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2039)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2039),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2040 transition  input  output  no-bypass 
    -- predecessors 500 
    -- successors 2041 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8255_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1701_base_resize_ack_0, ack => cp_elements(2040)); -- 
    sum_rename_req_8259_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2040), ack => ptr_deref_1701_root_address_inst_req_0); -- 
    -- CP-element group 2041 transition  input  output  no-bypass 
    -- predecessors 2040 
    -- successors 2042 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8260_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1701_root_address_inst_ack_0, ack => cp_elements(2041)); -- 
    root_register_req_8264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2041), ack => ptr_deref_1701_addr_0_req_0); -- 
    -- CP-element group 2042 fork  transition  input  no-bypass 
    -- predecessors 2041 
    -- successors 2038 2043 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_word_addrgen/root_register_ack
      -- 
    root_register_ack_8265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1701_addr_0_ack_0, ack => cp_elements(2042)); -- 
    -- CP-element group 2043 transition  output  bypass 
    -- predecessors 2042 
    -- successors 2044 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/word_access/word_access_0/rr
      -- 
    cp_elements(2043) <= cp_elements(2042);
    rr_8275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2043), ack => ptr_deref_1701_load_0_req_0); -- 
    -- CP-element group 2044 transition  input  no-bypass 
    -- predecessors 2043 
    -- successors 2038 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_request/word_access/word_access_0/ra
      -- 
    ra_8276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1701_load_0_ack_0, ack => cp_elements(2044)); -- 
    -- CP-element group 2045 transition  output  bypass 
    -- predecessors 2038 
    -- successors 2046 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2045) <= cp_elements(2038);
    cr_8286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2045), ack => ptr_deref_1701_load_0_req_1); -- 
    -- CP-element group 2046 transition  input  output  no-bypass 
    -- predecessors 2045 
    -- successors 2047 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/merge_req
      -- 
    ca_8287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1701_load_0_ack_1, ack => cp_elements(2046)); -- 
    merge_req_8288_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2046), ack => ptr_deref_1701_gather_scatter_req_0); -- 
    -- CP-element group 2047 transition  input  no-bypass 
    -- predecessors 2046 
    -- successors 2039 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1701_complete/merge_ack
      -- 
    merge_ack_8289_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1701_gather_scatter_ack_0, ack => cp_elements(2047)); -- 
    -- CP-element group 2048 join  fork  transition  bypass 
    -- predecessors 2052 2054 
    -- successors 2049 2055 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_active_
      -- 
    cpelement_group_2048 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2052);
      predecessors(1) <= cp_elements(2054);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2048)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2048),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2049 join  fork  transition  bypass 
    -- predecessors 2048 2057 
    -- successors 2096 2161 2226 2291 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1706_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1706_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1706_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_completed_
      -- 
    cpelement_group_2049 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2048);
      predecessors(1) <= cp_elements(2057);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2049)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2049),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2050 transition  input  output  no-bypass 
    -- predecessors 476 
    -- successors 2051 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1705_base_resize_ack_0, ack => cp_elements(2050)); -- 
    sum_rename_req_8311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2050), ack => ptr_deref_1705_root_address_inst_req_0); -- 
    -- CP-element group 2051 transition  input  output  no-bypass 
    -- predecessors 2050 
    -- successors 2052 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1705_root_address_inst_ack_0, ack => cp_elements(2051)); -- 
    root_register_req_8316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2051), ack => ptr_deref_1705_addr_0_req_0); -- 
    -- CP-element group 2052 fork  transition  input  no-bypass 
    -- predecessors 2051 
    -- successors 2048 2053 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_word_addrgen/root_register_ack
      -- 
    root_register_ack_8317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1705_addr_0_ack_0, ack => cp_elements(2052)); -- 
    -- CP-element group 2053 transition  output  bypass 
    -- predecessors 2052 
    -- successors 2054 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/word_access/word_access_0/rr
      -- 
    cp_elements(2053) <= cp_elements(2052);
    rr_8327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2053), ack => ptr_deref_1705_load_0_req_0); -- 
    -- CP-element group 2054 transition  input  no-bypass 
    -- predecessors 2053 
    -- successors 2048 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_request/word_access/word_access_0/ra
      -- 
    ra_8328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1705_load_0_ack_0, ack => cp_elements(2054)); -- 
    -- CP-element group 2055 transition  output  bypass 
    -- predecessors 2048 
    -- successors 2056 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2055) <= cp_elements(2048);
    cr_8338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2055), ack => ptr_deref_1705_load_0_req_1); -- 
    -- CP-element group 2056 transition  input  output  no-bypass 
    -- predecessors 2055 
    -- successors 2057 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/merge_req
      -- 
    ca_8339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1705_load_0_ack_1, ack => cp_elements(2056)); -- 
    merge_req_8340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2056), ack => ptr_deref_1705_gather_scatter_req_0); -- 
    -- CP-element group 2057 transition  input  no-bypass 
    -- predecessors 2056 
    -- successors 2049 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1705_complete/merge_ack
      -- 
    merge_ack_8341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1705_gather_scatter_ack_0, ack => cp_elements(2057)); -- 
    -- CP-element group 2058 join  fork  transition  bypass 
    -- predecessors 2062 2064 
    -- successors 2059 2065 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_active_
      -- 
    cpelement_group_2058 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2062);
      predecessors(1) <= cp_elements(2064);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2058)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2058),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2059 join  fork  transition  bypass 
    -- predecessors 2058 2067 
    -- successors 2105 2170 2235 2300 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1710_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1710_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1710_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_completed_
      -- 
    cpelement_group_2059 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2058);
      predecessors(1) <= cp_elements(2067);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2059)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2059),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2060 transition  input  output  no-bypass 
    -- predecessors 459 
    -- successors 2061 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1709_base_resize_ack_0, ack => cp_elements(2060)); -- 
    sum_rename_req_8363_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2060), ack => ptr_deref_1709_root_address_inst_req_0); -- 
    -- CP-element group 2061 transition  input  output  no-bypass 
    -- predecessors 2060 
    -- successors 2062 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8364_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1709_root_address_inst_ack_0, ack => cp_elements(2061)); -- 
    root_register_req_8368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2061), ack => ptr_deref_1709_addr_0_req_0); -- 
    -- CP-element group 2062 fork  transition  input  no-bypass 
    -- predecessors 2061 
    -- successors 2058 2063 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_word_addrgen/root_register_ack
      -- 
    root_register_ack_8369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1709_addr_0_ack_0, ack => cp_elements(2062)); -- 
    -- CP-element group 2063 transition  output  bypass 
    -- predecessors 2062 
    -- successors 2064 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/word_access/word_access_0/rr
      -- 
    cp_elements(2063) <= cp_elements(2062);
    rr_8379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2063), ack => ptr_deref_1709_load_0_req_0); -- 
    -- CP-element group 2064 transition  input  no-bypass 
    -- predecessors 2063 
    -- successors 2058 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_request/word_access/word_access_0/ra
      -- 
    ra_8380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1709_load_0_ack_0, ack => cp_elements(2064)); -- 
    -- CP-element group 2065 transition  output  bypass 
    -- predecessors 2058 
    -- successors 2066 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2065) <= cp_elements(2058);
    cr_8390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2065), ack => ptr_deref_1709_load_0_req_1); -- 
    -- CP-element group 2066 transition  input  output  no-bypass 
    -- predecessors 2065 
    -- successors 2067 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/merge_req
      -- 
    ca_8391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1709_load_0_ack_1, ack => cp_elements(2066)); -- 
    merge_req_8392_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2066), ack => ptr_deref_1709_gather_scatter_req_0); -- 
    -- CP-element group 2067 transition  input  no-bypass 
    -- predecessors 2066 
    -- successors 2059 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/ptr_deref_1709_complete/merge_ack
      -- 
    merge_ack_8393_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1709_gather_scatter_ack_0, ack => cp_elements(2067)); -- 
    -- CP-element group 2068 join  fork  transition  no-bypass 
    -- predecessors 2071 2072 
    -- successors 2069 2073 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_trigger_
      -- 
    cpelement_group_2068 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2071);
      predecessors(1) <= cp_elements(2072);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2068)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2068),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2069 join  fork  transition  no-bypass 
    -- predecessors 2068 2074 
    -- successors 2070 2075 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_active_
      -- 
    cpelement_group_2069 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2068);
      predecessors(1) <= cp_elements(2074);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2069)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2069),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2070 join  transition  bypass 
    -- predecessors 2069 2076 
    -- successors 2086 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1715_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1715_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1715_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1722_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1722_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1722_completed_
      -- 
    cpelement_group_2070 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2069);
      predecessors(1) <= cp_elements(2076);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2070)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2070),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2071 transition  bypass 
    -- predecessors 2029 
    -- successors 2068 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1712_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1712_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1712_completed_
      -- 
    cp_elements(2071) <= cp_elements(2029);
    -- CP-element group 2072 transition  bypass 
    -- predecessors 979 
    -- successors 2068 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1713_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1713_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1713_completed_
      -- 
    cp_elements(2072) <= cp_elements(979);
    -- CP-element group 2073 transition  output  bypass 
    -- predecessors 2068 
    -- successors 2074 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Sample/rr
      -- 
    cp_elements(2073) <= cp_elements(2068);
    rr_8409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2073), ack => binary_1714_inst_req_0); -- 
    -- CP-element group 2074 transition  input  no-bypass 
    -- predecessors 2073 
    -- successors 2069 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Sample/ra
      -- 
    ra_8410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1714_inst_ack_0, ack => cp_elements(2074)); -- 
    -- CP-element group 2075 transition  output  bypass 
    -- predecessors 2069 
    -- successors 2076 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Update/cr
      -- 
    cp_elements(2075) <= cp_elements(2069);
    cr_8414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2075), ack => binary_1714_inst_req_1); -- 
    -- CP-element group 2076 transition  input  no-bypass 
    -- predecessors 2075 
    -- successors 2070 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1714_complete_Update/ca
      -- 
    ca_8415_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1714_inst_ack_1, ack => cp_elements(2076)); -- 
    -- CP-element group 2077 join  fork  transition  no-bypass 
    -- predecessors 2080 2081 
    -- successors 2078 2082 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_trigger_
      -- 
    cpelement_group_2077 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2080);
      predecessors(1) <= cp_elements(2081);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2077)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2077),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2078 join  fork  transition  no-bypass 
    -- predecessors 2077 2083 
    -- successors 2079 2084 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_active_
      -- 
    cpelement_group_2078 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2077);
      predecessors(1) <= cp_elements(2083);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2078)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2078),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2079 join  transition  bypass 
    -- predecessors 2078 2085 
    -- successors 2086 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1720_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1720_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1720_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1723_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1723_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1723_completed_
      -- 
    cpelement_group_2079 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2078);
      predecessors(1) <= cp_elements(2085);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2079)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2079),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2080 transition  bypass 
    -- predecessors 2039 
    -- successors 2077 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1717_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1717_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1717_completed_
      -- 
    cp_elements(2080) <= cp_elements(2039);
    -- CP-element group 2081 transition  bypass 
    -- predecessors 999 
    -- successors 2077 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1718_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1718_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1718_completed_
      -- 
    cp_elements(2081) <= cp_elements(999);
    -- CP-element group 2082 transition  output  bypass 
    -- predecessors 2077 
    -- successors 2083 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Sample/rr
      -- 
    cp_elements(2082) <= cp_elements(2077);
    rr_8431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2082), ack => binary_1719_inst_req_0); -- 
    -- CP-element group 2083 transition  input  no-bypass 
    -- predecessors 2082 
    -- successors 2078 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Sample/ra
      -- 
    ra_8432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1719_inst_ack_0, ack => cp_elements(2083)); -- 
    -- CP-element group 2084 transition  output  bypass 
    -- predecessors 2078 
    -- successors 2085 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Update/cr
      -- 
    cp_elements(2084) <= cp_elements(2078);
    cr_8436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2084), ack => binary_1719_inst_req_1); -- 
    -- CP-element group 2085 transition  input  no-bypass 
    -- predecessors 2084 
    -- successors 2079 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1719_complete_Update/ca
      -- 
    ca_8437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1719_inst_ack_1, ack => cp_elements(2085)); -- 
    -- CP-element group 2086 join  fork  transition  bypass 
    -- predecessors 2070 2079 
    -- successors 2087 2089 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_trigger_
      -- 
    cpelement_group_2086 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2070);
      predecessors(1) <= cp_elements(2079);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2086)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2086),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2087 join  fork  transition  no-bypass 
    -- predecessors 2086 2090 
    -- successors 2088 2091 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_active_
      -- 
    cpelement_group_2087 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2086);
      predecessors(1) <= cp_elements(2090);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2087)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2087),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2088 join  transition  no-bypass 
    -- predecessors 2087 2092 
    -- successors 2118 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1725_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1725_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1725_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1742_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1742_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1742_completed_
      -- 
    cpelement_group_2088 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2087);
      predecessors(1) <= cp_elements(2092);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2088)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2088),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2089 transition  output  bypass 
    -- predecessors 2086 
    -- successors 2090 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Sample/rr
      -- 
    cp_elements(2089) <= cp_elements(2086);
    rr_8453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2089), ack => binary_1724_inst_req_0); -- 
    -- CP-element group 2090 transition  input  no-bypass 
    -- predecessors 2089 
    -- successors 2087 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Sample/ra
      -- 
    ra_8454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1724_inst_ack_0, ack => cp_elements(2090)); -- 
    -- CP-element group 2091 transition  output  bypass 
    -- predecessors 2087 
    -- successors 2092 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Update/cr
      -- 
    cp_elements(2091) <= cp_elements(2087);
    cr_8458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2091), ack => binary_1724_inst_req_1); -- 
    -- CP-element group 2092 transition  input  no-bypass 
    -- predecessors 2091 
    -- successors 2088 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1724_complete_Update/ca
      -- 
    ca_8459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1724_inst_ack_1, ack => cp_elements(2092)); -- 
    -- CP-element group 2093 join  fork  transition  no-bypass 
    -- predecessors 2096 2097 
    -- successors 2094 2098 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_trigger_
      -- 
    cpelement_group_2093 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2096);
      predecessors(1) <= cp_elements(2097);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2093)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2093),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2094 join  fork  transition  no-bypass 
    -- predecessors 2093 2099 
    -- successors 2095 2100 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_active_
      -- 
    cpelement_group_2094 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2093);
      predecessors(1) <= cp_elements(2099);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2094)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2094),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2095 join  transition  bypass 
    -- predecessors 2094 2101 
    -- successors 2111 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1730_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1730_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1730_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1737_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1737_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1737_completed_
      -- 
    cpelement_group_2095 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2094);
      predecessors(1) <= cp_elements(2101);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2095)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2095),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2096 transition  bypass 
    -- predecessors 2049 
    -- successors 2093 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1727_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1727_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1727_completed_
      -- 
    cp_elements(2096) <= cp_elements(2049);
    -- CP-element group 2097 transition  bypass 
    -- predecessors 1019 
    -- successors 2093 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1728_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1728_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1728_completed_
      -- 
    cp_elements(2097) <= cp_elements(1019);
    -- CP-element group 2098 transition  output  bypass 
    -- predecessors 2093 
    -- successors 2099 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Sample/rr
      -- 
    cp_elements(2098) <= cp_elements(2093);
    rr_8475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2098), ack => binary_1729_inst_req_0); -- 
    -- CP-element group 2099 transition  input  no-bypass 
    -- predecessors 2098 
    -- successors 2094 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Sample/ra
      -- 
    ra_8476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1729_inst_ack_0, ack => cp_elements(2099)); -- 
    -- CP-element group 2100 transition  output  bypass 
    -- predecessors 2094 
    -- successors 2101 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Update/cr
      -- 
    cp_elements(2100) <= cp_elements(2094);
    cr_8480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2100), ack => binary_1729_inst_req_1); -- 
    -- CP-element group 2101 transition  input  no-bypass 
    -- predecessors 2100 
    -- successors 2095 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1729_complete_Update/ca
      -- 
    ca_8481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1729_inst_ack_1, ack => cp_elements(2101)); -- 
    -- CP-element group 2102 join  fork  transition  no-bypass 
    -- predecessors 2105 2106 
    -- successors 2103 2107 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_trigger_
      -- 
    cpelement_group_2102 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2105);
      predecessors(1) <= cp_elements(2106);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2102)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2102),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2103 join  fork  transition  no-bypass 
    -- predecessors 2102 2108 
    -- successors 2104 2109 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_active_
      -- 
    cpelement_group_2103 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2102);
      predecessors(1) <= cp_elements(2108);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2103)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2104 join  transition  bypass 
    -- predecessors 2103 2110 
    -- successors 2111 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1735_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1735_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1735_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1738_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1738_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1738_completed_
      -- 
    cpelement_group_2104 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2103);
      predecessors(1) <= cp_elements(2110);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2104)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2104),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2105 transition  bypass 
    -- predecessors 2059 
    -- successors 2102 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1732_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1732_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1732_completed_
      -- 
    cp_elements(2105) <= cp_elements(2059);
    -- CP-element group 2106 transition  bypass 
    -- predecessors 1039 
    -- successors 2102 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1733_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1733_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1733_completed_
      -- 
    cp_elements(2106) <= cp_elements(1039);
    -- CP-element group 2107 transition  output  bypass 
    -- predecessors 2102 
    -- successors 2108 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Sample/rr
      -- 
    cp_elements(2107) <= cp_elements(2102);
    rr_8497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2107), ack => binary_1734_inst_req_0); -- 
    -- CP-element group 2108 transition  input  no-bypass 
    -- predecessors 2107 
    -- successors 2103 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Sample/ra
      -- 
    ra_8498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1734_inst_ack_0, ack => cp_elements(2108)); -- 
    -- CP-element group 2109 transition  output  bypass 
    -- predecessors 2103 
    -- successors 2110 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Update/cr
      -- 
    cp_elements(2109) <= cp_elements(2103);
    cr_8502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2109), ack => binary_1734_inst_req_1); -- 
    -- CP-element group 2110 transition  input  no-bypass 
    -- predecessors 2109 
    -- successors 2104 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1734_complete_Update/ca
      -- 
    ca_8503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1734_inst_ack_1, ack => cp_elements(2110)); -- 
    -- CP-element group 2111 join  fork  transition  bypass 
    -- predecessors 2095 2104 
    -- successors 2112 2114 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_trigger_
      -- 
    cpelement_group_2111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2095);
      predecessors(1) <= cp_elements(2104);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2111)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2112 join  fork  transition  no-bypass 
    -- predecessors 2111 2115 
    -- successors 2113 2116 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_active_
      -- 
    cpelement_group_2112 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2111);
      predecessors(1) <= cp_elements(2115);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2112)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2113 join  transition  no-bypass 
    -- predecessors 2112 2117 
    -- successors 2118 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1740_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1740_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1740_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1743_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1743_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1743_completed_
      -- 
    cpelement_group_2113 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2112);
      predecessors(1) <= cp_elements(2117);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2113)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2114 transition  output  bypass 
    -- predecessors 2111 
    -- successors 2115 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Sample/rr
      -- 
    cp_elements(2114) <= cp_elements(2111);
    rr_8519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2114), ack => binary_1739_inst_req_0); -- 
    -- CP-element group 2115 transition  input  no-bypass 
    -- predecessors 2114 
    -- successors 2112 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Sample/ra
      -- 
    ra_8520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1739_inst_ack_0, ack => cp_elements(2115)); -- 
    -- CP-element group 2116 transition  output  bypass 
    -- predecessors 2112 
    -- successors 2117 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Update/cr
      -- 
    cp_elements(2116) <= cp_elements(2112);
    cr_8524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2116), ack => binary_1739_inst_req_1); -- 
    -- CP-element group 2117 transition  input  no-bypass 
    -- predecessors 2116 
    -- successors 2113 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1739_complete_Update/ca
      -- 
    ca_8525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1739_inst_ack_1, ack => cp_elements(2117)); -- 
    -- CP-element group 2118 join  fork  transition  bypass 
    -- predecessors 2088 2113 
    -- successors 2119 2121 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_trigger_
      -- 
    cpelement_group_2118 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2088);
      predecessors(1) <= cp_elements(2113);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2118)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2119 join  fork  transition  no-bypass 
    -- predecessors 2118 2122 
    -- successors 2120 2123 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_active_
      -- 
    cpelement_group_2119 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2118);
      predecessors(1) <= cp_elements(2122);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2119)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2119),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2120 join  transition  no-bypass 
    -- predecessors 2119 2124 
    -- successors 2125 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1745_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1745_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1745_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1748_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1748_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1748_completed_
      -- 
    cpelement_group_2120 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2119);
      predecessors(1) <= cp_elements(2124);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2120)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2120),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2121 transition  output  bypass 
    -- predecessors 2118 
    -- successors 2122 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Sample/rr
      -- 
    cp_elements(2121) <= cp_elements(2118);
    rr_8541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2121), ack => binary_1744_inst_req_0); -- 
    -- CP-element group 2122 transition  input  no-bypass 
    -- predecessors 2121 
    -- successors 2119 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Sample/ra
      -- 
    ra_8542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1744_inst_ack_0, ack => cp_elements(2122)); -- 
    -- CP-element group 2123 transition  output  bypass 
    -- predecessors 2119 
    -- successors 2124 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Update/cr
      -- 
    cp_elements(2123) <= cp_elements(2119);
    cr_8546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2123), ack => binary_1744_inst_req_1); -- 
    -- CP-element group 2124 transition  input  no-bypass 
    -- predecessors 2123 
    -- successors 2120 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1744_complete_Update/ca
      -- 
    ca_8547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1744_inst_ack_1, ack => cp_elements(2124)); -- 
    -- CP-element group 2125 join  fork  transition  no-bypass 
    -- predecessors 2120 2128 
    -- successors 2126 2129 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_trigger_
      -- 
    cpelement_group_2125 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2120);
      predecessors(1) <= cp_elements(2128);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2125)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2125),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2126 join  fork  transition  bypass 
    -- predecessors 2125 2130 
    -- successors 2127 2131 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_active_
      -- 
    cpelement_group_2126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2125);
      predecessors(1) <= cp_elements(2130);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2126)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2127 join  transition  bypass 
    -- predecessors 2126 2132 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1750_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1750_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1750_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_completed_
      -- 
    cpelement_group_2127 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2126);
      predecessors(1) <= cp_elements(2132);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2127)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2127),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2128 transition  bypass 
    -- predecessors 367 
    -- successors 2125 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1747_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1747_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1747_completed_
      -- 
    cp_elements(2128) <= cp_elements(367);
    -- CP-element group 2129 transition  output  bypass 
    -- predecessors 2125 
    -- successors 2130 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Sample/rr
      -- 
    cp_elements(2129) <= cp_elements(2125);
    rr_8563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2129), ack => binary_1749_inst_req_0); -- 
    -- CP-element group 2130 transition  input  no-bypass 
    -- predecessors 2129 
    -- successors 2126 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Sample/ra
      -- 
    ra_8564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1749_inst_ack_0, ack => cp_elements(2130)); -- 
    -- CP-element group 2131 transition  output  bypass 
    -- predecessors 2126 
    -- successors 2132 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Update/cr
      -- 
    cp_elements(2131) <= cp_elements(2126);
    cr_8568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2131), ack => binary_1749_inst_req_1); -- 
    -- CP-element group 2132 transition  input  no-bypass 
    -- predecessors 2131 
    -- successors 2127 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1749_complete_Update/ca
      -- 
    ca_8569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1749_inst_ack_1, ack => cp_elements(2132)); -- 
    -- CP-element group 2133 join  fork  transition  no-bypass 
    -- predecessors 2136 2137 
    -- successors 2134 2138 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_trigger_
      -- 
    cpelement_group_2133 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2136);
      predecessors(1) <= cp_elements(2137);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2133)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2133),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2134 join  fork  transition  no-bypass 
    -- predecessors 2133 2139 
    -- successors 2135 2140 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_active_
      -- 
    cpelement_group_2134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2133);
      predecessors(1) <= cp_elements(2139);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2134)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2135 join  transition  bypass 
    -- predecessors 2134 2141 
    -- successors 2151 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1755_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1755_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1755_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1762_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1762_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1762_completed_
      -- 
    cpelement_group_2135 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2134);
      predecessors(1) <= cp_elements(2141);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2135)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2135),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2136 transition  bypass 
    -- predecessors 2029 
    -- successors 2133 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1752_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1752_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1752_completed_
      -- 
    cp_elements(2136) <= cp_elements(2029);
    -- CP-element group 2137 transition  bypass 
    -- predecessors 1114 
    -- successors 2133 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1753_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1753_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1753_completed_
      -- 
    cp_elements(2137) <= cp_elements(1114);
    -- CP-element group 2138 transition  output  bypass 
    -- predecessors 2133 
    -- successors 2139 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Sample/rr
      -- 
    cp_elements(2138) <= cp_elements(2133);
    rr_8585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2138), ack => binary_1754_inst_req_0); -- 
    -- CP-element group 2139 transition  input  no-bypass 
    -- predecessors 2138 
    -- successors 2134 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Sample/ra
      -- 
    ra_8586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1754_inst_ack_0, ack => cp_elements(2139)); -- 
    -- CP-element group 2140 transition  output  bypass 
    -- predecessors 2134 
    -- successors 2141 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Update/cr
      -- 
    cp_elements(2140) <= cp_elements(2134);
    cr_8590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2140), ack => binary_1754_inst_req_1); -- 
    -- CP-element group 2141 transition  input  no-bypass 
    -- predecessors 2140 
    -- successors 2135 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1754_complete_Update/ca
      -- 
    ca_8591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1754_inst_ack_1, ack => cp_elements(2141)); -- 
    -- CP-element group 2142 join  fork  transition  no-bypass 
    -- predecessors 2145 2146 
    -- successors 2143 2147 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_trigger_
      -- 
    cpelement_group_2142 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2145);
      predecessors(1) <= cp_elements(2146);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2142)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2142),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2143 join  fork  transition  no-bypass 
    -- predecessors 2142 2148 
    -- successors 2144 2149 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_active_
      -- 
    cpelement_group_2143 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2142);
      predecessors(1) <= cp_elements(2148);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2143)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2143),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2144 join  transition  bypass 
    -- predecessors 2143 2150 
    -- successors 2151 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1760_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1760_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1760_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1763_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1763_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1763_completed_
      -- 
    cpelement_group_2144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2143);
      predecessors(1) <= cp_elements(2150);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2144)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2145 transition  bypass 
    -- predecessors 2039 
    -- successors 2142 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1757_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1757_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1757_completed_
      -- 
    cp_elements(2145) <= cp_elements(2039);
    -- CP-element group 2146 transition  bypass 
    -- predecessors 1124 
    -- successors 2142 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1758_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1758_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1758_completed_
      -- 
    cp_elements(2146) <= cp_elements(1124);
    -- CP-element group 2147 transition  output  bypass 
    -- predecessors 2142 
    -- successors 2148 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Sample/rr
      -- 
    cp_elements(2147) <= cp_elements(2142);
    rr_8607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2147), ack => binary_1759_inst_req_0); -- 
    -- CP-element group 2148 transition  input  no-bypass 
    -- predecessors 2147 
    -- successors 2143 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Sample/ra
      -- 
    ra_8608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1759_inst_ack_0, ack => cp_elements(2148)); -- 
    -- CP-element group 2149 transition  output  bypass 
    -- predecessors 2143 
    -- successors 2150 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Update/cr
      -- 
    cp_elements(2149) <= cp_elements(2143);
    cr_8612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2149), ack => binary_1759_inst_req_1); -- 
    -- CP-element group 2150 transition  input  no-bypass 
    -- predecessors 2149 
    -- successors 2144 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1759_complete_Update/ca
      -- 
    ca_8613_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1759_inst_ack_1, ack => cp_elements(2150)); -- 
    -- CP-element group 2151 join  fork  transition  bypass 
    -- predecessors 2135 2144 
    -- successors 2152 2154 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_trigger_
      -- 
    cpelement_group_2151 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2135);
      predecessors(1) <= cp_elements(2144);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2151)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2151),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2152 join  fork  transition  no-bypass 
    -- predecessors 2151 2155 
    -- successors 2153 2156 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_active_
      -- 
    cpelement_group_2152 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2151);
      predecessors(1) <= cp_elements(2155);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2152)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2152),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2153 join  transition  no-bypass 
    -- predecessors 2152 2157 
    -- successors 2183 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1765_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1765_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1765_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1782_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1782_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1782_completed_
      -- 
    cpelement_group_2153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2152);
      predecessors(1) <= cp_elements(2157);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2153)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2154 transition  output  bypass 
    -- predecessors 2151 
    -- successors 2155 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Sample/rr
      -- 
    cp_elements(2154) <= cp_elements(2151);
    rr_8629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2154), ack => binary_1764_inst_req_0); -- 
    -- CP-element group 2155 transition  input  no-bypass 
    -- predecessors 2154 
    -- successors 2152 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Sample/ra
      -- 
    ra_8630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1764_inst_ack_0, ack => cp_elements(2155)); -- 
    -- CP-element group 2156 transition  output  bypass 
    -- predecessors 2152 
    -- successors 2157 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Update/cr
      -- 
    cp_elements(2156) <= cp_elements(2152);
    cr_8634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2156), ack => binary_1764_inst_req_1); -- 
    -- CP-element group 2157 transition  input  no-bypass 
    -- predecessors 2156 
    -- successors 2153 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1764_complete_Update/ca
      -- 
    ca_8635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1764_inst_ack_1, ack => cp_elements(2157)); -- 
    -- CP-element group 2158 join  fork  transition  no-bypass 
    -- predecessors 2161 2162 
    -- successors 2159 2163 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_trigger_
      -- 
    cpelement_group_2158 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2161);
      predecessors(1) <= cp_elements(2162);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2158)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2158),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2159 join  fork  transition  no-bypass 
    -- predecessors 2158 2164 
    -- successors 2160 2165 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_active_
      -- 
    cpelement_group_2159 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2158);
      predecessors(1) <= cp_elements(2164);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2159)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2159),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2160 join  transition  bypass 
    -- predecessors 2159 2166 
    -- successors 2176 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1770_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1770_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1770_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1777_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1777_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1777_completed_
      -- 
    cpelement_group_2160 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2159);
      predecessors(1) <= cp_elements(2166);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2160)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2161 transition  bypass 
    -- predecessors 2049 
    -- successors 2158 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1767_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1767_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1767_completed_
      -- 
    cp_elements(2161) <= cp_elements(2049);
    -- CP-element group 2162 transition  bypass 
    -- predecessors 1134 
    -- successors 2158 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1768_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1768_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1768_completed_
      -- 
    cp_elements(2162) <= cp_elements(1134);
    -- CP-element group 2163 transition  output  bypass 
    -- predecessors 2158 
    -- successors 2164 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Sample/rr
      -- 
    cp_elements(2163) <= cp_elements(2158);
    rr_8651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2163), ack => binary_1769_inst_req_0); -- 
    -- CP-element group 2164 transition  input  no-bypass 
    -- predecessors 2163 
    -- successors 2159 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Sample/ra
      -- 
    ra_8652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1769_inst_ack_0, ack => cp_elements(2164)); -- 
    -- CP-element group 2165 transition  output  bypass 
    -- predecessors 2159 
    -- successors 2166 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Update/cr
      -- 
    cp_elements(2165) <= cp_elements(2159);
    cr_8656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2165), ack => binary_1769_inst_req_1); -- 
    -- CP-element group 2166 transition  input  no-bypass 
    -- predecessors 2165 
    -- successors 2160 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1769_complete_Update/ca
      -- 
    ca_8657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1769_inst_ack_1, ack => cp_elements(2166)); -- 
    -- CP-element group 2167 join  fork  transition  no-bypass 
    -- predecessors 2170 2171 
    -- successors 2168 2172 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_trigger_
      -- 
    cpelement_group_2167 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2170);
      predecessors(1) <= cp_elements(2171);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2167)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2167),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2168 join  fork  transition  no-bypass 
    -- predecessors 2167 2173 
    -- successors 2169 2174 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_active_
      -- 
    cpelement_group_2168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2167);
      predecessors(1) <= cp_elements(2173);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2168)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2169 join  transition  bypass 
    -- predecessors 2168 2175 
    -- successors 2176 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1775_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1775_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1775_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1778_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1778_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1778_completed_
      -- 
    cpelement_group_2169 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2168);
      predecessors(1) <= cp_elements(2175);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2169)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2169),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2170 transition  bypass 
    -- predecessors 2059 
    -- successors 2167 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1772_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1772_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1772_completed_
      -- 
    cp_elements(2170) <= cp_elements(2059);
    -- CP-element group 2171 transition  bypass 
    -- predecessors 1144 
    -- successors 2167 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1773_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1773_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1773_completed_
      -- 
    cp_elements(2171) <= cp_elements(1144);
    -- CP-element group 2172 transition  output  bypass 
    -- predecessors 2167 
    -- successors 2173 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Sample/rr
      -- 
    cp_elements(2172) <= cp_elements(2167);
    rr_8673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2172), ack => binary_1774_inst_req_0); -- 
    -- CP-element group 2173 transition  input  no-bypass 
    -- predecessors 2172 
    -- successors 2168 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Sample/ra
      -- 
    ra_8674_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1774_inst_ack_0, ack => cp_elements(2173)); -- 
    -- CP-element group 2174 transition  output  bypass 
    -- predecessors 2168 
    -- successors 2175 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Update/cr
      -- 
    cp_elements(2174) <= cp_elements(2168);
    cr_8678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2174), ack => binary_1774_inst_req_1); -- 
    -- CP-element group 2175 transition  input  no-bypass 
    -- predecessors 2174 
    -- successors 2169 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1774_complete_Update/ca
      -- 
    ca_8679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1774_inst_ack_1, ack => cp_elements(2175)); -- 
    -- CP-element group 2176 join  fork  transition  bypass 
    -- predecessors 2160 2169 
    -- successors 2177 2179 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_trigger_
      -- 
    cpelement_group_2176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2160);
      predecessors(1) <= cp_elements(2169);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2176)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2177 join  fork  transition  no-bypass 
    -- predecessors 2176 2180 
    -- successors 2178 2181 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_active_
      -- 
    cpelement_group_2177 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2176);
      predecessors(1) <= cp_elements(2180);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2177)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2177),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2178 join  transition  no-bypass 
    -- predecessors 2177 2182 
    -- successors 2183 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1780_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1780_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1780_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1783_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1783_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1783_completed_
      -- 
    cpelement_group_2178 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2177);
      predecessors(1) <= cp_elements(2182);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2178)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2178),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2179 transition  output  bypass 
    -- predecessors 2176 
    -- successors 2180 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Sample/rr
      -- 
    cp_elements(2179) <= cp_elements(2176);
    rr_8695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2179), ack => binary_1779_inst_req_0); -- 
    -- CP-element group 2180 transition  input  no-bypass 
    -- predecessors 2179 
    -- successors 2177 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Sample/ra
      -- 
    ra_8696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1779_inst_ack_0, ack => cp_elements(2180)); -- 
    -- CP-element group 2181 transition  output  bypass 
    -- predecessors 2177 
    -- successors 2182 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Update/cr
      -- 
    cp_elements(2181) <= cp_elements(2177);
    cr_8700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2181), ack => binary_1779_inst_req_1); -- 
    -- CP-element group 2182 transition  input  no-bypass 
    -- predecessors 2181 
    -- successors 2178 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1779_complete_Update/ca
      -- 
    ca_8701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1779_inst_ack_1, ack => cp_elements(2182)); -- 
    -- CP-element group 2183 join  fork  transition  bypass 
    -- predecessors 2153 2178 
    -- successors 2184 2186 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_trigger_
      -- 
    cpelement_group_2183 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2153);
      predecessors(1) <= cp_elements(2178);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2183)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2183),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2184 join  fork  transition  no-bypass 
    -- predecessors 2183 2187 
    -- successors 2185 2188 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_active_
      -- 
    cpelement_group_2184 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2183);
      predecessors(1) <= cp_elements(2187);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2184)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2184),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2185 join  transition  no-bypass 
    -- predecessors 2184 2189 
    -- successors 2190 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1785_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1785_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1785_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1788_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1788_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1788_completed_
      -- 
    cpelement_group_2185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2184);
      predecessors(1) <= cp_elements(2189);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2185)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2186 transition  output  bypass 
    -- predecessors 2183 
    -- successors 2187 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Sample/rr
      -- 
    cp_elements(2186) <= cp_elements(2183);
    rr_8717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2186), ack => binary_1784_inst_req_0); -- 
    -- CP-element group 2187 transition  input  no-bypass 
    -- predecessors 2186 
    -- successors 2184 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Sample/ra
      -- 
    ra_8718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1784_inst_ack_0, ack => cp_elements(2187)); -- 
    -- CP-element group 2188 transition  output  bypass 
    -- predecessors 2184 
    -- successors 2189 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Update/cr
      -- 
    cp_elements(2188) <= cp_elements(2184);
    cr_8722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2188), ack => binary_1784_inst_req_1); -- 
    -- CP-element group 2189 transition  input  no-bypass 
    -- predecessors 2188 
    -- successors 2185 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1784_complete_Update/ca
      -- 
    ca_8723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1784_inst_ack_1, ack => cp_elements(2189)); -- 
    -- CP-element group 2190 join  fork  transition  no-bypass 
    -- predecessors 2185 2193 
    -- successors 2191 2194 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_trigger_
      -- 
    cpelement_group_2190 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2185);
      predecessors(1) <= cp_elements(2193);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2190)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2190),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2191 join  fork  transition  bypass 
    -- predecessors 2190 2195 
    -- successors 2192 2196 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_active_
      -- 
    cpelement_group_2191 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2190);
      predecessors(1) <= cp_elements(2195);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2191)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2191),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2192 join  transition  bypass 
    -- predecessors 2191 2197 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1790_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1790_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1790_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_completed_
      -- 
    cpelement_group_2192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2191);
      predecessors(1) <= cp_elements(2197);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2192)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2193 transition  bypass 
    -- predecessors 367 
    -- successors 2190 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1787_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1787_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1787_completed_
      -- 
    cp_elements(2193) <= cp_elements(367);
    -- CP-element group 2194 transition  output  bypass 
    -- predecessors 2190 
    -- successors 2195 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Sample/rr
      -- 
    cp_elements(2194) <= cp_elements(2190);
    rr_8739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2194), ack => binary_1789_inst_req_0); -- 
    -- CP-element group 2195 transition  input  no-bypass 
    -- predecessors 2194 
    -- successors 2191 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Sample/ra
      -- 
    ra_8740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1789_inst_ack_0, ack => cp_elements(2195)); -- 
    -- CP-element group 2196 transition  output  bypass 
    -- predecessors 2191 
    -- successors 2197 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Update/cr
      -- 
    cp_elements(2196) <= cp_elements(2191);
    cr_8744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2196), ack => binary_1789_inst_req_1); -- 
    -- CP-element group 2197 transition  input  no-bypass 
    -- predecessors 2196 
    -- successors 2192 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1789_complete_Update/ca
      -- 
    ca_8745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1789_inst_ack_1, ack => cp_elements(2197)); -- 
    -- CP-element group 2198 join  fork  transition  no-bypass 
    -- predecessors 2201 2202 
    -- successors 2199 2203 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_trigger_
      -- 
    cpelement_group_2198 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2201);
      predecessors(1) <= cp_elements(2202);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2198)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2198),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2199 join  fork  transition  no-bypass 
    -- predecessors 2198 2204 
    -- successors 2200 2205 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_active_
      -- 
    cpelement_group_2199 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2198);
      predecessors(1) <= cp_elements(2204);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2199)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2200 join  transition  bypass 
    -- predecessors 2199 2206 
    -- successors 2216 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1802_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1802_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1802_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1795_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1795_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1795_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_completed_
      -- 
    cpelement_group_2200 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2199);
      predecessors(1) <= cp_elements(2206);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2200)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2200),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2201 transition  bypass 
    -- predecessors 2029 
    -- successors 2198 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1792_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1792_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1792_completed_
      -- 
    cp_elements(2201) <= cp_elements(2029);
    -- CP-element group 2202 transition  bypass 
    -- predecessors 1219 
    -- successors 2198 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1793_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1793_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1793_completed_
      -- 
    cp_elements(2202) <= cp_elements(1219);
    -- CP-element group 2203 transition  output  bypass 
    -- predecessors 2198 
    -- successors 2204 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Sample/rr
      -- 
    cp_elements(2203) <= cp_elements(2198);
    rr_8761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2203), ack => binary_1794_inst_req_0); -- 
    -- CP-element group 2204 transition  input  no-bypass 
    -- predecessors 2203 
    -- successors 2199 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Sample/ra
      -- 
    ra_8762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1794_inst_ack_0, ack => cp_elements(2204)); -- 
    -- CP-element group 2205 transition  output  bypass 
    -- predecessors 2199 
    -- successors 2206 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Update/cr
      -- 
    cp_elements(2205) <= cp_elements(2199);
    cr_8766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2205), ack => binary_1794_inst_req_1); -- 
    -- CP-element group 2206 transition  input  no-bypass 
    -- predecessors 2205 
    -- successors 2200 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1794_complete_Update/ca
      -- 
    ca_8767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1794_inst_ack_1, ack => cp_elements(2206)); -- 
    -- CP-element group 2207 join  fork  transition  no-bypass 
    -- predecessors 2210 2211 
    -- successors 2208 2212 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_trigger_
      -- 
    cpelement_group_2207 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2210);
      predecessors(1) <= cp_elements(2211);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2207)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2207),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2208 join  fork  transition  no-bypass 
    -- predecessors 2207 2213 
    -- successors 2209 2214 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_active_
      -- 
    cpelement_group_2208 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2207);
      predecessors(1) <= cp_elements(2213);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2208)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2208),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2209 join  transition  bypass 
    -- predecessors 2208 2215 
    -- successors 2216 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1803_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1803_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1803_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1800_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1800_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1800_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_completed_
      -- 
    cpelement_group_2209 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2208);
      predecessors(1) <= cp_elements(2215);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2209)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2209),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2210 transition  bypass 
    -- predecessors 2039 
    -- successors 2207 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1797_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1797_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1797_completed_
      -- 
    cp_elements(2210) <= cp_elements(2039);
    -- CP-element group 2211 transition  bypass 
    -- predecessors 1229 
    -- successors 2207 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1798_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1798_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1798_completed_
      -- 
    cp_elements(2211) <= cp_elements(1229);
    -- CP-element group 2212 transition  output  bypass 
    -- predecessors 2207 
    -- successors 2213 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Sample/rr
      -- 
    cp_elements(2212) <= cp_elements(2207);
    rr_8783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2212), ack => binary_1799_inst_req_0); -- 
    -- CP-element group 2213 transition  input  no-bypass 
    -- predecessors 2212 
    -- successors 2208 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Sample/ra
      -- 
    ra_8784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1799_inst_ack_0, ack => cp_elements(2213)); -- 
    -- CP-element group 2214 transition  output  bypass 
    -- predecessors 2208 
    -- successors 2215 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Update/cr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Update/$entry
      -- 
    cp_elements(2214) <= cp_elements(2208);
    cr_8788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2214), ack => binary_1799_inst_req_1); -- 
    -- CP-element group 2215 transition  input  no-bypass 
    -- predecessors 2214 
    -- successors 2209 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Update/ca
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1799_complete_Update/$exit
      -- 
    ca_8789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1799_inst_ack_1, ack => cp_elements(2215)); -- 
    -- CP-element group 2216 join  fork  transition  bypass 
    -- predecessors 2200 2209 
    -- successors 2217 2219 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_trigger_
      -- 
    cpelement_group_2216 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2200);
      predecessors(1) <= cp_elements(2209);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2216)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2216),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2217 join  fork  transition  no-bypass 
    -- predecessors 2216 2220 
    -- successors 2218 2221 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_active_
      -- 
    cpelement_group_2217 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2216);
      predecessors(1) <= cp_elements(2220);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2217)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2217),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2218 join  transition  no-bypass 
    -- predecessors 2217 2222 
    -- successors 2248 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1805_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1805_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1805_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1822_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1822_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1822_completed_
      -- 
    cpelement_group_2218 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2217);
      predecessors(1) <= cp_elements(2222);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2218)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2218),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2219 transition  output  bypass 
    -- predecessors 2216 
    -- successors 2220 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Sample/rr
      -- 
    cp_elements(2219) <= cp_elements(2216);
    rr_8805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2219), ack => binary_1804_inst_req_0); -- 
    -- CP-element group 2220 transition  input  no-bypass 
    -- predecessors 2219 
    -- successors 2217 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Sample/ra
      -- 
    ra_8806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1804_inst_ack_0, ack => cp_elements(2220)); -- 
    -- CP-element group 2221 transition  output  bypass 
    -- predecessors 2217 
    -- successors 2222 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Update/cr
      -- 
    cp_elements(2221) <= cp_elements(2217);
    cr_8810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2221), ack => binary_1804_inst_req_1); -- 
    -- CP-element group 2222 transition  input  no-bypass 
    -- predecessors 2221 
    -- successors 2218 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1804_complete_Update/ca
      -- 
    ca_8811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1804_inst_ack_1, ack => cp_elements(2222)); -- 
    -- CP-element group 2223 join  fork  transition  no-bypass 
    -- predecessors 2226 2227 
    -- successors 2224 2228 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_trigger_
      -- 
    cpelement_group_2223 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2226);
      predecessors(1) <= cp_elements(2227);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2223)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2223),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2224 join  fork  transition  no-bypass 
    -- predecessors 2223 2229 
    -- successors 2225 2230 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_active_
      -- 
    cpelement_group_2224 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2223);
      predecessors(1) <= cp_elements(2229);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2224)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2224),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2225 join  transition  bypass 
    -- predecessors 2224 2231 
    -- successors 2241 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1817_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1817_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1810_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1810_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1810_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1817_completed_
      -- 
    cpelement_group_2225 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2224);
      predecessors(1) <= cp_elements(2231);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2225)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2225),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2226 transition  bypass 
    -- predecessors 2049 
    -- successors 2223 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1807_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1807_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1807_completed_
      -- 
    cp_elements(2226) <= cp_elements(2049);
    -- CP-element group 2227 transition  bypass 
    -- predecessors 1239 
    -- successors 2223 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1808_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1808_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1808_completed_
      -- 
    cp_elements(2227) <= cp_elements(1239);
    -- CP-element group 2228 transition  output  bypass 
    -- predecessors 2223 
    -- successors 2229 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Sample/rr
      -- 
    cp_elements(2228) <= cp_elements(2223);
    rr_8827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2228), ack => binary_1809_inst_req_0); -- 
    -- CP-element group 2229 transition  input  no-bypass 
    -- predecessors 2228 
    -- successors 2224 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Sample/ra
      -- 
    ra_8828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1809_inst_ack_0, ack => cp_elements(2229)); -- 
    -- CP-element group 2230 transition  output  bypass 
    -- predecessors 2224 
    -- successors 2231 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Update/cr
      -- 
    cp_elements(2230) <= cp_elements(2224);
    cr_8832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2230), ack => binary_1809_inst_req_1); -- 
    -- CP-element group 2231 transition  input  no-bypass 
    -- predecessors 2230 
    -- successors 2225 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1809_complete_Update/ca
      -- 
    ca_8833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1809_inst_ack_1, ack => cp_elements(2231)); -- 
    -- CP-element group 2232 join  fork  transition  no-bypass 
    -- predecessors 2235 2236 
    -- successors 2233 2237 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_trigger_
      -- 
    cpelement_group_2232 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2235);
      predecessors(1) <= cp_elements(2236);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2232)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2232),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2233 join  fork  transition  no-bypass 
    -- predecessors 2232 2238 
    -- successors 2234 2239 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_active_
      -- 
    cpelement_group_2233 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2232);
      predecessors(1) <= cp_elements(2238);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2233)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2233),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2234 join  transition  bypass 
    -- predecessors 2233 2240 
    -- successors 2241 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1818_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1818_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1815_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1815_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1815_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1818_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_completed_
      -- 
    cpelement_group_2234 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2233);
      predecessors(1) <= cp_elements(2240);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2234)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2234),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2235 transition  bypass 
    -- predecessors 2059 
    -- successors 2232 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1812_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1812_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1812_trigger_
      -- 
    cp_elements(2235) <= cp_elements(2059);
    -- CP-element group 2236 transition  bypass 
    -- predecessors 1249 
    -- successors 2232 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1813_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1813_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1813_completed_
      -- 
    cp_elements(2236) <= cp_elements(1249);
    -- CP-element group 2237 transition  output  bypass 
    -- predecessors 2232 
    -- successors 2238 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Sample/rr
      -- 
    cp_elements(2237) <= cp_elements(2232);
    rr_8849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2237), ack => binary_1814_inst_req_0); -- 
    -- CP-element group 2238 transition  input  no-bypass 
    -- predecessors 2237 
    -- successors 2233 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Sample/ra
      -- 
    ra_8850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1814_inst_ack_0, ack => cp_elements(2238)); -- 
    -- CP-element group 2239 transition  output  bypass 
    -- predecessors 2233 
    -- successors 2240 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Update/cr
      -- 
    cp_elements(2239) <= cp_elements(2233);
    cr_8854_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2239), ack => binary_1814_inst_req_1); -- 
    -- CP-element group 2240 transition  input  no-bypass 
    -- predecessors 2239 
    -- successors 2234 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1814_complete_Update/ca
      -- 
    ca_8855_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1814_inst_ack_1, ack => cp_elements(2240)); -- 
    -- CP-element group 2241 join  fork  transition  bypass 
    -- predecessors 2225 2234 
    -- successors 2242 2244 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_trigger_
      -- 
    cpelement_group_2241 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2225);
      predecessors(1) <= cp_elements(2234);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2241)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2241),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2242 join  fork  transition  no-bypass 
    -- predecessors 2241 2245 
    -- successors 2243 2246 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_active_
      -- 
    cpelement_group_2242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2241);
      predecessors(1) <= cp_elements(2245);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2242)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2243 join  transition  no-bypass 
    -- predecessors 2242 2247 
    -- successors 2248 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1820_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1820_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1820_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1823_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1823_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1823_completed_
      -- 
    cpelement_group_2243 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2242);
      predecessors(1) <= cp_elements(2247);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2243)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2243),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2244 transition  output  bypass 
    -- predecessors 2241 
    -- successors 2245 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Sample/rr
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Sample/$entry
      -- 
    cp_elements(2244) <= cp_elements(2241);
    rr_8871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2244), ack => binary_1819_inst_req_0); -- 
    -- CP-element group 2245 transition  input  no-bypass 
    -- predecessors 2244 
    -- successors 2242 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Sample/ra
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Sample/$exit
      -- 
    ra_8872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1819_inst_ack_0, ack => cp_elements(2245)); -- 
    -- CP-element group 2246 transition  output  bypass 
    -- predecessors 2242 
    -- successors 2247 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Update/cr
      -- 
    cp_elements(2246) <= cp_elements(2242);
    cr_8876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2246), ack => binary_1819_inst_req_1); -- 
    -- CP-element group 2247 transition  input  no-bypass 
    -- predecessors 2246 
    -- successors 2243 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1819_complete_Update/ca
      -- 
    ca_8877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1819_inst_ack_1, ack => cp_elements(2247)); -- 
    -- CP-element group 2248 join  fork  transition  bypass 
    -- predecessors 2218 2243 
    -- successors 2249 2251 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_trigger_
      -- 
    cpelement_group_2248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2218);
      predecessors(1) <= cp_elements(2243);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2248)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2249 join  fork  transition  no-bypass 
    -- predecessors 2248 2252 
    -- successors 2250 2253 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_active_
      -- 
    cpelement_group_2249 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2248);
      predecessors(1) <= cp_elements(2252);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2249)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2249),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2250 join  transition  no-bypass 
    -- predecessors 2249 2254 
    -- successors 2255 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1825_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1825_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1825_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1828_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1828_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1828_completed_
      -- 
    cpelement_group_2250 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2249);
      predecessors(1) <= cp_elements(2254);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2250)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2250),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2251 transition  output  bypass 
    -- predecessors 2248 
    -- successors 2252 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Sample/rr
      -- 
    cp_elements(2251) <= cp_elements(2248);
    rr_8893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2251), ack => binary_1824_inst_req_0); -- 
    -- CP-element group 2252 transition  input  no-bypass 
    -- predecessors 2251 
    -- successors 2249 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Sample/ra
      -- 
    ra_8894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1824_inst_ack_0, ack => cp_elements(2252)); -- 
    -- CP-element group 2253 transition  output  bypass 
    -- predecessors 2249 
    -- successors 2254 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Update/cr
      -- 
    cp_elements(2253) <= cp_elements(2249);
    cr_8898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2253), ack => binary_1824_inst_req_1); -- 
    -- CP-element group 2254 transition  input  no-bypass 
    -- predecessors 2253 
    -- successors 2250 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1824_complete_Update/ca
      -- 
    ca_8899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1824_inst_ack_1, ack => cp_elements(2254)); -- 
    -- CP-element group 2255 join  fork  transition  no-bypass 
    -- predecessors 2250 2258 
    -- successors 2256 2259 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_trigger_
      -- 
    cpelement_group_2255 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2250);
      predecessors(1) <= cp_elements(2258);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2255)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2256 join  fork  transition  bypass 
    -- predecessors 2255 2260 
    -- successors 2257 2261 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_active_
      -- 
    cpelement_group_2256 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2255);
      predecessors(1) <= cp_elements(2260);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2256)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2256),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2257 join  transition  bypass 
    -- predecessors 2256 2262 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1830_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1830_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1830_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_completed_
      -- 
    cpelement_group_2257 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2256);
      predecessors(1) <= cp_elements(2262);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2257)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2257),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2258 transition  bypass 
    -- predecessors 367 
    -- successors 2255 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1827_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1827_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1827_completed_
      -- 
    cp_elements(2258) <= cp_elements(367);
    -- CP-element group 2259 transition  output  bypass 
    -- predecessors 2255 
    -- successors 2260 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Sample/rr
      -- 
    cp_elements(2259) <= cp_elements(2255);
    rr_8915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2259), ack => binary_1829_inst_req_0); -- 
    -- CP-element group 2260 transition  input  no-bypass 
    -- predecessors 2259 
    -- successors 2256 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Sample/ra
      -- 
    ra_8916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1829_inst_ack_0, ack => cp_elements(2260)); -- 
    -- CP-element group 2261 transition  output  bypass 
    -- predecessors 2256 
    -- successors 2262 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Update/cr
      -- 
    cp_elements(2261) <= cp_elements(2256);
    cr_8920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2261), ack => binary_1829_inst_req_1); -- 
    -- CP-element group 2262 transition  input  no-bypass 
    -- predecessors 2261 
    -- successors 2257 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1829_complete_Update/ca
      -- 
    ca_8921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1829_inst_ack_1, ack => cp_elements(2262)); -- 
    -- CP-element group 2263 join  fork  transition  no-bypass 
    -- predecessors 2266 2267 
    -- successors 2264 2268 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_trigger_
      -- 
    cpelement_group_2263 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2266);
      predecessors(1) <= cp_elements(2267);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2263)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2263),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2264 join  fork  transition  no-bypass 
    -- predecessors 2263 2269 
    -- successors 2265 2270 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_active_
      -- 
    cpelement_group_2264 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2263);
      predecessors(1) <= cp_elements(2269);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2264)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2264),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2265 join  transition  bypass 
    -- predecessors 2264 2271 
    -- successors 2281 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1835_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1835_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1835_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1842_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1842_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1842_completed_
      -- 
    cpelement_group_2265 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2264);
      predecessors(1) <= cp_elements(2271);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2265)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2265),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2266 transition  bypass 
    -- predecessors 2029 
    -- successors 2263 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1832_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1832_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1832_completed_
      -- 
    cp_elements(2266) <= cp_elements(2029);
    -- CP-element group 2267 transition  bypass 
    -- predecessors 1324 
    -- successors 2263 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1833_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1833_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1833_completed_
      -- 
    cp_elements(2267) <= cp_elements(1324);
    -- CP-element group 2268 transition  output  bypass 
    -- predecessors 2263 
    -- successors 2269 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Sample/rr
      -- 
    cp_elements(2268) <= cp_elements(2263);
    rr_8937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2268), ack => binary_1834_inst_req_0); -- 
    -- CP-element group 2269 transition  input  no-bypass 
    -- predecessors 2268 
    -- successors 2264 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Sample/ra
      -- 
    ra_8938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1834_inst_ack_0, ack => cp_elements(2269)); -- 
    -- CP-element group 2270 transition  output  bypass 
    -- predecessors 2264 
    -- successors 2271 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Update/cr
      -- 
    cp_elements(2270) <= cp_elements(2264);
    cr_8942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2270), ack => binary_1834_inst_req_1); -- 
    -- CP-element group 2271 transition  input  no-bypass 
    -- predecessors 2270 
    -- successors 2265 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1834_complete_Update/ca
      -- 
    ca_8943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1834_inst_ack_1, ack => cp_elements(2271)); -- 
    -- CP-element group 2272 join  fork  transition  no-bypass 
    -- predecessors 2275 2276 
    -- successors 2273 2277 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_trigger_
      -- 
    cpelement_group_2272 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2275);
      predecessors(1) <= cp_elements(2276);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2272)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2273 join  fork  transition  no-bypass 
    -- predecessors 2272 2278 
    -- successors 2274 2279 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_active_
      -- 
    cpelement_group_2273 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2272);
      predecessors(1) <= cp_elements(2278);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2273)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2273),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2274 join  transition  bypass 
    -- predecessors 2273 2280 
    -- successors 2281 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1840_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1840_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1840_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1843_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1843_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1843_completed_
      -- 
    cpelement_group_2274 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2273);
      predecessors(1) <= cp_elements(2280);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2274)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2274),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2275 transition  bypass 
    -- predecessors 2039 
    -- successors 2272 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1837_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1837_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1837_completed_
      -- 
    cp_elements(2275) <= cp_elements(2039);
    -- CP-element group 2276 transition  bypass 
    -- predecessors 1334 
    -- successors 2272 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1838_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1838_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1838_completed_
      -- 
    cp_elements(2276) <= cp_elements(1334);
    -- CP-element group 2277 transition  output  bypass 
    -- predecessors 2272 
    -- successors 2278 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Sample/rr
      -- 
    cp_elements(2277) <= cp_elements(2272);
    rr_8959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2277), ack => binary_1839_inst_req_0); -- 
    -- CP-element group 2278 transition  input  no-bypass 
    -- predecessors 2277 
    -- successors 2273 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Sample/ra
      -- 
    ra_8960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1839_inst_ack_0, ack => cp_elements(2278)); -- 
    -- CP-element group 2279 transition  output  bypass 
    -- predecessors 2273 
    -- successors 2280 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Update/cr
      -- 
    cp_elements(2279) <= cp_elements(2273);
    cr_8964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2279), ack => binary_1839_inst_req_1); -- 
    -- CP-element group 2280 transition  input  no-bypass 
    -- predecessors 2279 
    -- successors 2274 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1839_complete_Update/ca
      -- 
    ca_8965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1839_inst_ack_1, ack => cp_elements(2280)); -- 
    -- CP-element group 2281 join  fork  transition  bypass 
    -- predecessors 2265 2274 
    -- successors 2282 2284 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_trigger_
      -- 
    cpelement_group_2281 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2265);
      predecessors(1) <= cp_elements(2274);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2281)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2282 join  fork  transition  no-bypass 
    -- predecessors 2281 2285 
    -- successors 2283 2286 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_active_
      -- 
    cpelement_group_2282 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2281);
      predecessors(1) <= cp_elements(2285);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2282)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2282),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2283 join  transition  no-bypass 
    -- predecessors 2282 2287 
    -- successors 2313 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1845_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1845_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1845_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1862_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1862_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1862_completed_
      -- 
    cpelement_group_2283 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2282);
      predecessors(1) <= cp_elements(2287);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2283)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2283),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2284 transition  output  bypass 
    -- predecessors 2281 
    -- successors 2285 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Sample/rr
      -- 
    cp_elements(2284) <= cp_elements(2281);
    rr_8981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2284), ack => binary_1844_inst_req_0); -- 
    -- CP-element group 2285 transition  input  no-bypass 
    -- predecessors 2284 
    -- successors 2282 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Sample/ra
      -- 
    ra_8982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1844_inst_ack_0, ack => cp_elements(2285)); -- 
    -- CP-element group 2286 transition  output  bypass 
    -- predecessors 2282 
    -- successors 2287 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Update/cr
      -- 
    cp_elements(2286) <= cp_elements(2282);
    cr_8986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2286), ack => binary_1844_inst_req_1); -- 
    -- CP-element group 2287 transition  input  no-bypass 
    -- predecessors 2286 
    -- successors 2283 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1844_complete_Update/ca
      -- 
    ca_8987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1844_inst_ack_1, ack => cp_elements(2287)); -- 
    -- CP-element group 2288 join  fork  transition  no-bypass 
    -- predecessors 2291 2292 
    -- successors 2289 2293 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_trigger_
      -- 
    cpelement_group_2288 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2291);
      predecessors(1) <= cp_elements(2292);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2288)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2288),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2289 join  fork  transition  no-bypass 
    -- predecessors 2288 2294 
    -- successors 2290 2295 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_active_
      -- 
    cpelement_group_2289 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2288);
      predecessors(1) <= cp_elements(2294);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2289)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2289),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2290 join  transition  bypass 
    -- predecessors 2289 2296 
    -- successors 2306 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1850_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1850_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1850_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1857_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1857_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1857_completed_
      -- 
    cpelement_group_2290 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2289);
      predecessors(1) <= cp_elements(2296);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2290)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2291 transition  bypass 
    -- predecessors 2049 
    -- successors 2288 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1847_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1847_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1847_completed_
      -- 
    cp_elements(2291) <= cp_elements(2049);
    -- CP-element group 2292 transition  bypass 
    -- predecessors 1344 
    -- successors 2288 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1848_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1848_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1848_completed_
      -- 
    cp_elements(2292) <= cp_elements(1344);
    -- CP-element group 2293 transition  output  bypass 
    -- predecessors 2288 
    -- successors 2294 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Sample/rr
      -- 
    cp_elements(2293) <= cp_elements(2288);
    rr_9003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2293), ack => binary_1849_inst_req_0); -- 
    -- CP-element group 2294 transition  input  no-bypass 
    -- predecessors 2293 
    -- successors 2289 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Sample/ra
      -- 
    ra_9004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1849_inst_ack_0, ack => cp_elements(2294)); -- 
    -- CP-element group 2295 transition  output  bypass 
    -- predecessors 2289 
    -- successors 2296 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Update/cr
      -- 
    cp_elements(2295) <= cp_elements(2289);
    cr_9008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2295), ack => binary_1849_inst_req_1); -- 
    -- CP-element group 2296 transition  input  no-bypass 
    -- predecessors 2295 
    -- successors 2290 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1849_complete_Update/ca
      -- 
    ca_9009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1849_inst_ack_1, ack => cp_elements(2296)); -- 
    -- CP-element group 2297 join  fork  transition  no-bypass 
    -- predecessors 2300 2301 
    -- successors 2298 2302 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_trigger_
      -- 
    cpelement_group_2297 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2300);
      predecessors(1) <= cp_elements(2301);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2297)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2297),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2298 join  fork  transition  no-bypass 
    -- predecessors 2297 2303 
    -- successors 2299 2304 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_active_
      -- 
    cpelement_group_2298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2297);
      predecessors(1) <= cp_elements(2303);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2298)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2299 join  transition  bypass 
    -- predecessors 2298 2305 
    -- successors 2306 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1855_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1855_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1855_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1858_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1858_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1858_completed_
      -- 
    cpelement_group_2299 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2298);
      predecessors(1) <= cp_elements(2305);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2299)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2299),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2300 transition  bypass 
    -- predecessors 2059 
    -- successors 2297 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1852_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1852_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1852_completed_
      -- 
    cp_elements(2300) <= cp_elements(2059);
    -- CP-element group 2301 transition  bypass 
    -- predecessors 1354 
    -- successors 2297 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1853_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1853_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1853_completed_
      -- 
    cp_elements(2301) <= cp_elements(1354);
    -- CP-element group 2302 transition  output  bypass 
    -- predecessors 2297 
    -- successors 2303 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Sample/rr
      -- 
    cp_elements(2302) <= cp_elements(2297);
    rr_9025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2302), ack => binary_1854_inst_req_0); -- 
    -- CP-element group 2303 transition  input  no-bypass 
    -- predecessors 2302 
    -- successors 2298 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Sample/ra
      -- 
    ra_9026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1854_inst_ack_0, ack => cp_elements(2303)); -- 
    -- CP-element group 2304 transition  output  bypass 
    -- predecessors 2298 
    -- successors 2305 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Update/cr
      -- 
    cp_elements(2304) <= cp_elements(2298);
    cr_9030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2304), ack => binary_1854_inst_req_1); -- 
    -- CP-element group 2305 transition  input  no-bypass 
    -- predecessors 2304 
    -- successors 2299 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1854_complete_Update/ca
      -- 
    ca_9031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1854_inst_ack_1, ack => cp_elements(2305)); -- 
    -- CP-element group 2306 join  fork  transition  bypass 
    -- predecessors 2290 2299 
    -- successors 2307 2309 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_trigger_
      -- 
    cpelement_group_2306 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2290);
      predecessors(1) <= cp_elements(2299);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2306)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2306),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2307 join  fork  transition  no-bypass 
    -- predecessors 2306 2310 
    -- successors 2308 2311 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_active_
      -- 
    cpelement_group_2307 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2306);
      predecessors(1) <= cp_elements(2310);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2307)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2307),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2308 join  transition  no-bypass 
    -- predecessors 2307 2312 
    -- successors 2313 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1860_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1860_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1860_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1863_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1863_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1863_completed_
      -- 
    cpelement_group_2308 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2307);
      predecessors(1) <= cp_elements(2312);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2308)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2309 transition  output  bypass 
    -- predecessors 2306 
    -- successors 2310 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Sample/rr
      -- 
    cp_elements(2309) <= cp_elements(2306);
    rr_9047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2309), ack => binary_1859_inst_req_0); -- 
    -- CP-element group 2310 transition  input  no-bypass 
    -- predecessors 2309 
    -- successors 2307 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Sample/ra
      -- 
    ra_9048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1859_inst_ack_0, ack => cp_elements(2310)); -- 
    -- CP-element group 2311 transition  output  bypass 
    -- predecessors 2307 
    -- successors 2312 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Update/cr
      -- 
    cp_elements(2311) <= cp_elements(2307);
    cr_9052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2311), ack => binary_1859_inst_req_1); -- 
    -- CP-element group 2312 transition  input  no-bypass 
    -- predecessors 2311 
    -- successors 2308 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1859_complete_Update/ca
      -- 
    ca_9053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1859_inst_ack_1, ack => cp_elements(2312)); -- 
    -- CP-element group 2313 join  fork  transition  bypass 
    -- predecessors 2283 2308 
    -- successors 2314 2316 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_trigger_
      -- 
    cpelement_group_2313 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2283);
      predecessors(1) <= cp_elements(2308);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2313)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2313),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2314 join  fork  transition  no-bypass 
    -- predecessors 2313 2317 
    -- successors 2315 2318 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_active_
      -- 
    cpelement_group_2314 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2313);
      predecessors(1) <= cp_elements(2317);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2314)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2314),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2315 join  transition  no-bypass 
    -- predecessors 2314 2319 
    -- successors 2320 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1865_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1865_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1865_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1868_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1868_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1868_completed_
      -- 
    cpelement_group_2315 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2314);
      predecessors(1) <= cp_elements(2319);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2315)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2315),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2316 transition  output  bypass 
    -- predecessors 2313 
    -- successors 2317 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Sample/rr
      -- 
    cp_elements(2316) <= cp_elements(2313);
    rr_9069_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2316), ack => binary_1864_inst_req_0); -- 
    -- CP-element group 2317 transition  input  no-bypass 
    -- predecessors 2316 
    -- successors 2314 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Sample/ra
      -- 
    ra_9070_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1864_inst_ack_0, ack => cp_elements(2317)); -- 
    -- CP-element group 2318 transition  output  bypass 
    -- predecessors 2314 
    -- successors 2319 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Update/cr
      -- 
    cp_elements(2318) <= cp_elements(2314);
    cr_9074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2318), ack => binary_1864_inst_req_1); -- 
    -- CP-element group 2319 transition  input  no-bypass 
    -- predecessors 2318 
    -- successors 2315 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1864_complete_Update/ca
      -- 
    ca_9075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1864_inst_ack_1, ack => cp_elements(2319)); -- 
    -- CP-element group 2320 join  fork  transition  no-bypass 
    -- predecessors 2315 2323 
    -- successors 2321 2324 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_trigger_
      -- 
    cpelement_group_2320 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2315);
      predecessors(1) <= cp_elements(2323);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2320)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2320),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2321 join  fork  transition  bypass 
    -- predecessors 2320 2325 
    -- successors 2322 2326 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_active_
      -- 
    cpelement_group_2321 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2320);
      predecessors(1) <= cp_elements(2325);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2321)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2321),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2322 join  transition  bypass 
    -- predecessors 2321 2327 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1870_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1870_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1870_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_completed_
      -- 
    cpelement_group_2322 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2321);
      predecessors(1) <= cp_elements(2327);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2322)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2322),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2323 transition  bypass 
    -- predecessors 367 
    -- successors 2320 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1867_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1867_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1867_completed_
      -- 
    cp_elements(2323) <= cp_elements(367);
    -- CP-element group 2324 transition  output  bypass 
    -- predecessors 2320 
    -- successors 2325 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Sample/rr
      -- 
    cp_elements(2324) <= cp_elements(2320);
    rr_9091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2324), ack => binary_1869_inst_req_0); -- 
    -- CP-element group 2325 transition  input  no-bypass 
    -- predecessors 2324 
    -- successors 2321 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Sample/ra
      -- 
    ra_9092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1869_inst_ack_0, ack => cp_elements(2325)); -- 
    -- CP-element group 2326 transition  output  bypass 
    -- predecessors 2321 
    -- successors 2327 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Update/cr
      -- 
    cp_elements(2326) <= cp_elements(2321);
    cr_9096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2326), ack => binary_1869_inst_req_1); -- 
    -- CP-element group 2327 transition  input  no-bypass 
    -- predecessors 2326 
    -- successors 2322 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1869_complete_Update/ca
      -- 
    ca_9097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1869_inst_ack_1, ack => cp_elements(2327)); -- 
    -- CP-element group 2328 join  fork  transition  no-bypass 
    -- predecessors 2330 2332 
    -- successors 2329 2333 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_active_
      -- 
    cpelement_group_2328 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2330);
      predecessors(1) <= cp_elements(2332);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2328)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2328),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2329 join  fork  transition  bypass 
    -- predecessors 2328 2334 
    -- successors 2335 2337 
    -- members (8) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1876_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1876_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1876_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1878_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1878_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1878_completed_
      -- 
    cpelement_group_2329 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2328);
      predecessors(1) <= cp_elements(2334);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2329)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2329),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2330 fork  transition  bypass 
    -- predecessors 367 
    -- successors 2328 2331 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1872_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1872_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/simple_obj_ref_1872_completed_
      -- 
    cp_elements(2330) <= cp_elements(367);
    -- CP-element group 2331 transition  output  bypass 
    -- predecessors 2330 
    -- successors 2332 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Sample/rr
      -- 
    cp_elements(2331) <= cp_elements(2330);
    rr_9110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2331), ack => binary_1875_inst_req_0); -- 
    -- CP-element group 2332 transition  input  no-bypass 
    -- predecessors 2331 
    -- successors 2328 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Sample/ra
      -- 
    ra_9111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1875_inst_ack_0, ack => cp_elements(2332)); -- 
    -- CP-element group 2333 transition  output  bypass 
    -- predecessors 2328 
    -- successors 2334 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Update/cr
      -- 
    cp_elements(2333) <= cp_elements(2328);
    cr_9115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2333), ack => binary_1875_inst_req_1); -- 
    -- CP-element group 2334 transition  input  no-bypass 
    -- predecessors 2333 
    -- successors 2329 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1875_complete_Update/ca
      -- 
    ca_9116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1875_inst_ack_1, ack => cp_elements(2334)); -- 
    -- CP-element group 2335 join  fork  transition  bypass 
    -- predecessors 2329 2338 
    -- successors 2336 2339 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_active_
      -- 
    cpelement_group_2335 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2329);
      predecessors(1) <= cp_elements(2338);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2335)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2335),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2336 join  transition  no-bypass 
    -- predecessors 2335 2340 
    -- successors 2341 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1882_trigger_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1882_active_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/assign_stmt_1882_completed_
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_completed_
      -- 
    cpelement_group_2336 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2335);
      predecessors(1) <= cp_elements(2340);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2336)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2336),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2337 transition  output  bypass 
    -- predecessors 2329 
    -- successors 2338 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Sample/rr
      -- 
    cp_elements(2337) <= cp_elements(2329);
    rr_9129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2337), ack => binary_1881_inst_req_0); -- 
    -- CP-element group 2338 transition  input  no-bypass 
    -- predecessors 2337 
    -- successors 2335 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Sample/ra
      -- 
    ra_9130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1881_inst_ack_0, ack => cp_elements(2338)); -- 
    -- CP-element group 2339 transition  output  bypass 
    -- predecessors 2335 
    -- successors 2340 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Update/cr
      -- 
    cp_elements(2339) <= cp_elements(2335);
    cr_9134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2339), ack => binary_1881_inst_req_1); -- 
    -- CP-element group 2340 transition  input  no-bypass 
    -- predecessors 2339 
    -- successors 2336 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/binary_1881_complete_Update/ca
      -- 
    ca_9135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1881_inst_ack_1, ack => cp_elements(2340)); -- 
    -- CP-element group 2341 join  transition  no-bypass 
    -- predecessors 1107 1212 1317 1422 1527 1592 1657 1722 1827 1892 1957 2022 2127 2192 2257 2322 2336 
    -- successors 4 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_868_to_assign_stmt_1882/$exit
      -- 
    cpelement_group_2341 : Block -- 
      signal predecessors: BooleanArray(16 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1107);
      predecessors(1) <= cp_elements(1212);
      predecessors(2) <= cp_elements(1317);
      predecessors(3) <= cp_elements(1422);
      predecessors(4) <= cp_elements(1527);
      predecessors(5) <= cp_elements(1592);
      predecessors(6) <= cp_elements(1657);
      predecessors(7) <= cp_elements(1722);
      predecessors(8) <= cp_elements(1827);
      predecessors(9) <= cp_elements(1892);
      predecessors(10) <= cp_elements(1957);
      predecessors(11) <= cp_elements(2022);
      predecessors(12) <= cp_elements(2127);
      predecessors(13) <= cp_elements(2192);
      predecessors(14) <= cp_elements(2257);
      predecessors(15) <= cp_elements(2322);
      predecessors(16) <= cp_elements(2336);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2341)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2341),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2342 transition  bypass 
    -- predecessors 4 
    -- successors 2343 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_1883_dead_link/$entry
      -- 
    cp_elements(2342) <= cp_elements(4);
    -- CP-element group 2343 transition  dead  bypass 
    -- predecessors 2342 
    -- successors 2344 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_1883_dead_link/dead_transition
      -- 
    cp_elements(2343) <= false;
    -- CP-element group 2344 transition  place  bypass 
    -- predecessors 2343 
    -- successors 2719 
    -- members (4) 
      -- 	branch_block_stmt_552/merge_stmt_1889__entry__
      -- 	branch_block_stmt_552/if_stmt_1883__exit__
      -- 	branch_block_stmt_552/if_stmt_1883_dead_link/$exit
      -- 	branch_block_stmt_552/merge_stmt_1889_dead_link/$entry
      -- 
    cp_elements(2344) <= cp_elements(2343);
    -- CP-element group 2345 transition  output  bypass 
    -- predecessors 4 
    -- successors 2346 
    -- members (3) 
      -- 	branch_block_stmt_552/if_stmt_1883_eval_test/$entry
      -- 	branch_block_stmt_552/if_stmt_1883_eval_test/$exit
      -- 	branch_block_stmt_552/if_stmt_1883_eval_test/branch_req
      -- 
    cp_elements(2345) <= cp_elements(4);
    branch_req_9143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2345), ack => if_stmt_1883_branch_req_0); -- 
    -- CP-element group 2346 branch  place  bypass 
    -- predecessors 2345 
    -- successors 2347 2349 
    -- members (1) 
      -- 	branch_block_stmt_552/simple_obj_ref_1884_place
      -- 
    cp_elements(2346) <= cp_elements(2345);
    -- CP-element group 2347 transition  bypass 
    -- predecessors 2346 
    -- successors 2348 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_1883_if_link/$entry
      -- 
    cp_elements(2347) <= cp_elements(2346);
    -- CP-element group 2348 transition  place  input  no-bypass 
    -- predecessors 2347 
    -- successors 2721 
    -- members (3) 
      -- 	branch_block_stmt_552/if_stmt_1883_if_link/$exit
      -- 	branch_block_stmt_552/if_stmt_1883_if_link/if_choice_transition
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge
      -- 
    if_choice_transition_9148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1883_branch_ack_1, ack => cp_elements(2348)); -- 
    -- CP-element group 2349 transition  bypass 
    -- predecessors 2346 
    -- successors 2350 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_1883_else_link/$entry
      -- 
    cp_elements(2349) <= cp_elements(2346);
    -- CP-element group 2350 transition  place  input  no-bypass 
    -- predecessors 2349 
    -- successors 2644 
    -- members (3) 
      -- 	branch_block_stmt_552/if_stmt_1883_else_link/$exit
      -- 	branch_block_stmt_552/if_stmt_1883_else_link/else_choice_transition
      -- 	branch_block_stmt_552/bb_3_bb_3
      -- 
    else_choice_transition_9152_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1883_branch_ack_0, ack => cp_elements(2350)); -- 
    -- CP-element group 2351 fork  transition  bypass 
    -- predecessors 5 
    -- successors 2353 2357 2368 2372 2383 2387 2398 2402 2413 2417 2428 2432 2443 2447 2458 2462 2473 2477 2488 2492 2503 2507 2518 2522 2533 2537 2548 2552 2563 2567 2578 2582 2594 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/$entry
      -- 
    cp_elements(2351) <= cp_elements(5);
    -- CP-element group 2352 join  transition  no-bypass 
    -- predecessors 2353 2356 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1958_completed_
      -- 
    cpelement_group_2352 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2353);
      predecessors(1) <= cp_elements(2356);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2352)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2352),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2353 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2352 2354 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1958_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1958_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1957_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1957_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1957_completed_
      -- 
    cp_elements(2353) <= cp_elements(2351);
    -- CP-element group 2354 join  fork  transition  no-bypass 
    -- predecessors 2353 2357 2361 
    -- successors 2355 2362 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_trigger_
      -- 
    cpelement_group_2354 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2353);
      predecessors(1) <= cp_elements(2357);
      predecessors(2) <= cp_elements(2361);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2354)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2354),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2355 join  fork  transition  bypass 
    -- predecessors 2354 2364 
    -- successors 2356 2365 2369 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_active_
      -- 
    cpelement_group_2355 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2354);
      predecessors(1) <= cp_elements(2364);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2355)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2355),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2356 join  transition  bypass 
    -- predecessors 2355 2366 
    -- successors 2352 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_completed_
      -- 
    cpelement_group_2356 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2355);
      predecessors(1) <= cp_elements(2366);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2356)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2356),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2357 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2354 2358 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1955_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1955_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1955_completed_
      -- 
    cp_elements(2357) <= cp_elements(2351);
    -- CP-element group 2358 transition  output  bypass 
    -- predecessors 2357 
    -- successors 2359 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_addr_resize/base_resize_req
      -- 
    cp_elements(2358) <= cp_elements(2357);
    base_resize_req_9177_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2358), ack => ptr_deref_1956_base_resize_req_0); -- 
    -- CP-element group 2359 transition  input  output  no-bypass 
    -- predecessors 2358 
    -- successors 2360 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1956_base_resize_ack_0, ack => cp_elements(2359)); -- 
    sum_rename_req_9182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2359), ack => ptr_deref_1956_root_address_inst_req_0); -- 
    -- CP-element group 2360 transition  input  output  no-bypass 
    -- predecessors 2359 
    -- successors 2361 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1956_root_address_inst_ack_0, ack => cp_elements(2360)); -- 
    root_register_req_9187_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2360), ack => ptr_deref_1956_addr_0_req_0); -- 
    -- CP-element group 2361 transition  input  no-bypass 
    -- predecessors 2360 
    -- successors 2354 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_word_addrgen/root_register_ack
      -- 
    root_register_ack_9188_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1956_addr_0_ack_0, ack => cp_elements(2361)); -- 
    -- CP-element group 2362 transition  output  bypass 
    -- predecessors 2354 
    -- successors 2363 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/split_req
      -- 
    cp_elements(2362) <= cp_elements(2354);
    split_req_9192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2362), ack => ptr_deref_1956_gather_scatter_req_0); -- 
    -- CP-element group 2363 transition  input  output  no-bypass 
    -- predecessors 2362 
    -- successors 2364 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/word_access/word_access_0/rr
      -- 
    split_ack_9193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1956_gather_scatter_ack_0, ack => cp_elements(2363)); -- 
    rr_9200_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2363), ack => ptr_deref_1956_store_0_req_0); -- 
    -- CP-element group 2364 transition  input  no-bypass 
    -- predecessors 2363 
    -- successors 2355 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_request/word_access/word_access_0/ra
      -- 
    ra_9201_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1956_store_0_ack_0, ack => cp_elements(2364)); -- 
    -- CP-element group 2365 transition  output  bypass 
    -- predecessors 2355 
    -- successors 2366 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2365) <= cp_elements(2355);
    cr_9211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2365), ack => ptr_deref_1956_store_0_req_1); -- 
    -- CP-element group 2366 transition  input  no-bypass 
    -- predecessors 2365 
    -- successors 2356 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1956_complete/word_access/word_access_0/ca
      -- 
    ca_9212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1956_store_0_ack_1, ack => cp_elements(2366)); -- 
    -- CP-element group 2367 join  transition  no-bypass 
    -- predecessors 2368 2371 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1962_completed_
      -- 
    cpelement_group_2367 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2368);
      predecessors(1) <= cp_elements(2371);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2367)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2367),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2368 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2367 2369 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1962_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1962_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1961_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1961_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1961_completed_
      -- 
    cp_elements(2368) <= cp_elements(2351);
    -- CP-element group 2369 join  fork  transition  no-bypass 
    -- predecessors 2355 2368 2372 2376 
    -- successors 2370 2377 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_trigger_
      -- 
    cpelement_group_2369 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2355);
      predecessors(1) <= cp_elements(2368);
      predecessors(2) <= cp_elements(2372);
      predecessors(3) <= cp_elements(2376);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2369)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2369),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2370 join  fork  transition  bypass 
    -- predecessors 2369 2379 
    -- successors 2371 2380 2384 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_active_
      -- 
    cpelement_group_2370 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2369);
      predecessors(1) <= cp_elements(2379);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2370)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2370),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2371 join  transition  bypass 
    -- predecessors 2370 2381 
    -- successors 2367 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_completed_
      -- 
    cpelement_group_2371 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2370);
      predecessors(1) <= cp_elements(2381);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2371)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2371),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2372 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2369 2373 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1959_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1959_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1959_completed_
      -- 
    cp_elements(2372) <= cp_elements(2351);
    -- CP-element group 2373 transition  output  bypass 
    -- predecessors 2372 
    -- successors 2374 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_addr_resize/base_resize_req
      -- 
    cp_elements(2373) <= cp_elements(2372);
    base_resize_req_9232_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2373), ack => ptr_deref_1960_base_resize_req_0); -- 
    -- CP-element group 2374 transition  input  output  no-bypass 
    -- predecessors 2373 
    -- successors 2375 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9233_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1960_base_resize_ack_0, ack => cp_elements(2374)); -- 
    sum_rename_req_9237_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2374), ack => ptr_deref_1960_root_address_inst_req_0); -- 
    -- CP-element group 2375 transition  input  output  no-bypass 
    -- predecessors 2374 
    -- successors 2376 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1960_root_address_inst_ack_0, ack => cp_elements(2375)); -- 
    root_register_req_9242_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2375), ack => ptr_deref_1960_addr_0_req_0); -- 
    -- CP-element group 2376 transition  input  no-bypass 
    -- predecessors 2375 
    -- successors 2369 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_word_addrgen/root_register_ack
      -- 
    root_register_ack_9243_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1960_addr_0_ack_0, ack => cp_elements(2376)); -- 
    -- CP-element group 2377 transition  output  bypass 
    -- predecessors 2369 
    -- successors 2378 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/split_req
      -- 
    cp_elements(2377) <= cp_elements(2369);
    split_req_9247_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2377), ack => ptr_deref_1960_gather_scatter_req_0); -- 
    -- CP-element group 2378 transition  input  output  no-bypass 
    -- predecessors 2377 
    -- successors 2379 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/word_access/word_access_0/rr
      -- 
    split_ack_9248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1960_gather_scatter_ack_0, ack => cp_elements(2378)); -- 
    rr_9255_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2378), ack => ptr_deref_1960_store_0_req_0); -- 
    -- CP-element group 2379 transition  input  no-bypass 
    -- predecessors 2378 
    -- successors 2370 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_request/word_access/word_access_0/ra
      -- 
    ra_9256_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1960_store_0_ack_0, ack => cp_elements(2379)); -- 
    -- CP-element group 2380 transition  output  bypass 
    -- predecessors 2370 
    -- successors 2381 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2380) <= cp_elements(2370);
    cr_9266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2380), ack => ptr_deref_1960_store_0_req_1); -- 
    -- CP-element group 2381 transition  input  no-bypass 
    -- predecessors 2380 
    -- successors 2371 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1960_complete/word_access/word_access_0/ca
      -- 
    ca_9267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1960_store_0_ack_1, ack => cp_elements(2381)); -- 
    -- CP-element group 2382 join  transition  no-bypass 
    -- predecessors 2383 2386 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1966_completed_
      -- 
    cpelement_group_2382 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2383);
      predecessors(1) <= cp_elements(2386);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2382)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2382),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2383 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2382 2384 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1966_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1966_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1965_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1965_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1965_completed_
      -- 
    cp_elements(2383) <= cp_elements(2351);
    -- CP-element group 2384 join  fork  transition  no-bypass 
    -- predecessors 2370 2383 2387 2391 
    -- successors 2385 2392 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_trigger_
      -- 
    cpelement_group_2384 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2370);
      predecessors(1) <= cp_elements(2383);
      predecessors(2) <= cp_elements(2387);
      predecessors(3) <= cp_elements(2391);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2384)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2384),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2385 join  fork  transition  bypass 
    -- predecessors 2384 2394 
    -- successors 2386 2395 2399 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_active_
      -- 
    cpelement_group_2385 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2384);
      predecessors(1) <= cp_elements(2394);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2385)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2385),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2386 join  transition  bypass 
    -- predecessors 2385 2396 
    -- successors 2382 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_completed_
      -- 
    cpelement_group_2386 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2385);
      predecessors(1) <= cp_elements(2396);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2386)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2386),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2387 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2384 2388 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1963_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1963_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1963_completed_
      -- 
    cp_elements(2387) <= cp_elements(2351);
    -- CP-element group 2388 transition  output  bypass 
    -- predecessors 2387 
    -- successors 2389 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_addr_resize/base_resize_req
      -- 
    cp_elements(2388) <= cp_elements(2387);
    base_resize_req_9287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2388), ack => ptr_deref_1964_base_resize_req_0); -- 
    -- CP-element group 2389 transition  input  output  no-bypass 
    -- predecessors 2388 
    -- successors 2390 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9288_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_base_resize_ack_0, ack => cp_elements(2389)); -- 
    sum_rename_req_9292_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2389), ack => ptr_deref_1964_root_address_inst_req_0); -- 
    -- CP-element group 2390 transition  input  output  no-bypass 
    -- predecessors 2389 
    -- successors 2391 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9293_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_root_address_inst_ack_0, ack => cp_elements(2390)); -- 
    root_register_req_9297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2390), ack => ptr_deref_1964_addr_0_req_0); -- 
    -- CP-element group 2391 transition  input  no-bypass 
    -- predecessors 2390 
    -- successors 2384 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_word_addrgen/root_register_ack
      -- 
    root_register_ack_9298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_addr_0_ack_0, ack => cp_elements(2391)); -- 
    -- CP-element group 2392 transition  output  bypass 
    -- predecessors 2384 
    -- successors 2393 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/split_req
      -- 
    cp_elements(2392) <= cp_elements(2384);
    split_req_9302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2392), ack => ptr_deref_1964_gather_scatter_req_0); -- 
    -- CP-element group 2393 transition  input  output  no-bypass 
    -- predecessors 2392 
    -- successors 2394 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/word_access/word_access_0/rr
      -- 
    split_ack_9303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_gather_scatter_ack_0, ack => cp_elements(2393)); -- 
    rr_9310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2393), ack => ptr_deref_1964_store_0_req_0); -- 
    -- CP-element group 2394 transition  input  no-bypass 
    -- predecessors 2393 
    -- successors 2385 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_request/word_access/word_access_0/ra
      -- 
    ra_9311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_store_0_ack_0, ack => cp_elements(2394)); -- 
    -- CP-element group 2395 transition  output  bypass 
    -- predecessors 2385 
    -- successors 2396 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2395) <= cp_elements(2385);
    cr_9321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2395), ack => ptr_deref_1964_store_0_req_1); -- 
    -- CP-element group 2396 transition  input  no-bypass 
    -- predecessors 2395 
    -- successors 2386 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1964_complete/word_access/word_access_0/ca
      -- 
    ca_9322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1964_store_0_ack_1, ack => cp_elements(2396)); -- 
    -- CP-element group 2397 join  transition  no-bypass 
    -- predecessors 2398 2401 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1970_completed_
      -- 
    cpelement_group_2397 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2398);
      predecessors(1) <= cp_elements(2401);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2397)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2397),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2398 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2397 2399 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1969_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1969_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1969_completed_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1970_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1970_active_
      -- 
    cp_elements(2398) <= cp_elements(2351);
    -- CP-element group 2399 join  fork  transition  no-bypass 
    -- predecessors 2385 2398 2402 2406 
    -- successors 2400 2407 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_trigger_
      -- 
    cpelement_group_2399 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2385);
      predecessors(1) <= cp_elements(2398);
      predecessors(2) <= cp_elements(2402);
      predecessors(3) <= cp_elements(2406);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2399)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2399),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2400 join  fork  transition  bypass 
    -- predecessors 2399 2409 
    -- successors 2401 2410 2414 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_active_
      -- 
    cpelement_group_2400 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2399);
      predecessors(1) <= cp_elements(2409);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2400)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2400),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2401 join  transition  bypass 
    -- predecessors 2400 2411 
    -- successors 2397 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_completed_
      -- 
    cpelement_group_2401 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2400);
      predecessors(1) <= cp_elements(2411);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2401)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2401),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2402 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2399 2403 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1967_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1967_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1967_completed_
      -- 
    cp_elements(2402) <= cp_elements(2351);
    -- CP-element group 2403 transition  output  bypass 
    -- predecessors 2402 
    -- successors 2404 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_addr_resize/base_resize_req
      -- 
    cp_elements(2403) <= cp_elements(2402);
    base_resize_req_9342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2403), ack => ptr_deref_1968_base_resize_req_0); -- 
    -- CP-element group 2404 transition  input  output  no-bypass 
    -- predecessors 2403 
    -- successors 2405 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_base_resize_ack_0, ack => cp_elements(2404)); -- 
    sum_rename_req_9347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2404), ack => ptr_deref_1968_root_address_inst_req_0); -- 
    -- CP-element group 2405 transition  input  output  no-bypass 
    -- predecessors 2404 
    -- successors 2406 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_root_address_inst_ack_0, ack => cp_elements(2405)); -- 
    root_register_req_9352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2405), ack => ptr_deref_1968_addr_0_req_0); -- 
    -- CP-element group 2406 transition  input  no-bypass 
    -- predecessors 2405 
    -- successors 2399 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_word_addrgen/root_register_ack
      -- 
    root_register_ack_9353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_addr_0_ack_0, ack => cp_elements(2406)); -- 
    -- CP-element group 2407 transition  output  bypass 
    -- predecessors 2399 
    -- successors 2408 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/split_req
      -- 
    cp_elements(2407) <= cp_elements(2399);
    split_req_9357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2407), ack => ptr_deref_1968_gather_scatter_req_0); -- 
    -- CP-element group 2408 transition  input  output  no-bypass 
    -- predecessors 2407 
    -- successors 2409 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/word_access/word_access_0/rr
      -- 
    split_ack_9358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_gather_scatter_ack_0, ack => cp_elements(2408)); -- 
    rr_9365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2408), ack => ptr_deref_1968_store_0_req_0); -- 
    -- CP-element group 2409 transition  input  no-bypass 
    -- predecessors 2408 
    -- successors 2400 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_request/word_access/word_access_0/ra
      -- 
    ra_9366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_store_0_ack_0, ack => cp_elements(2409)); -- 
    -- CP-element group 2410 transition  output  bypass 
    -- predecessors 2400 
    -- successors 2411 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2410) <= cp_elements(2400);
    cr_9376_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2410), ack => ptr_deref_1968_store_0_req_1); -- 
    -- CP-element group 2411 transition  input  no-bypass 
    -- predecessors 2410 
    -- successors 2401 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1968_complete/word_access/word_access_0/ca
      -- 
    ca_9377_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1968_store_0_ack_1, ack => cp_elements(2411)); -- 
    -- CP-element group 2412 join  transition  no-bypass 
    -- predecessors 2413 2416 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1974_completed_
      -- 
    cpelement_group_2412 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2413);
      predecessors(1) <= cp_elements(2416);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2412)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2412),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2413 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2412 2414 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1974_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1974_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1973_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1973_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1973_completed_
      -- 
    cp_elements(2413) <= cp_elements(2351);
    -- CP-element group 2414 join  fork  transition  no-bypass 
    -- predecessors 2400 2413 2417 2421 
    -- successors 2415 2422 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_trigger_
      -- 
    cpelement_group_2414 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2400);
      predecessors(1) <= cp_elements(2413);
      predecessors(2) <= cp_elements(2417);
      predecessors(3) <= cp_elements(2421);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2414)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2414),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2415 join  fork  transition  bypass 
    -- predecessors 2414 2424 
    -- successors 2416 2425 2429 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_active_
      -- 
    cpelement_group_2415 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2414);
      predecessors(1) <= cp_elements(2424);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2415)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2415),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2416 join  transition  bypass 
    -- predecessors 2415 2426 
    -- successors 2412 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_completed_
      -- 
    cpelement_group_2416 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2415);
      predecessors(1) <= cp_elements(2426);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2416)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2416),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2417 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2414 2418 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1971_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1971_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1971_completed_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_address_calculated
      -- 
    cp_elements(2417) <= cp_elements(2351);
    -- CP-element group 2418 transition  output  bypass 
    -- predecessors 2417 
    -- successors 2419 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_addr_resize/base_resize_req
      -- 
    cp_elements(2418) <= cp_elements(2417);
    base_resize_req_9397_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2418), ack => ptr_deref_1972_base_resize_req_0); -- 
    -- CP-element group 2419 transition  input  output  no-bypass 
    -- predecessors 2418 
    -- successors 2420 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9398_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_base_resize_ack_0, ack => cp_elements(2419)); -- 
    sum_rename_req_9402_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2419), ack => ptr_deref_1972_root_address_inst_req_0); -- 
    -- CP-element group 2420 transition  input  output  no-bypass 
    -- predecessors 2419 
    -- successors 2421 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9403_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_root_address_inst_ack_0, ack => cp_elements(2420)); -- 
    root_register_req_9407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2420), ack => ptr_deref_1972_addr_0_req_0); -- 
    -- CP-element group 2421 transition  input  no-bypass 
    -- predecessors 2420 
    -- successors 2414 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_word_addrgen/root_register_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_word_address_calculated
      -- 
    root_register_ack_9408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_0_ack_0, ack => cp_elements(2421)); -- 
    -- CP-element group 2422 transition  output  bypass 
    -- predecessors 2414 
    -- successors 2423 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/split_req
      -- 
    cp_elements(2422) <= cp_elements(2414);
    split_req_9412_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2422), ack => ptr_deref_1972_gather_scatter_req_0); -- 
    -- CP-element group 2423 transition  input  output  no-bypass 
    -- predecessors 2422 
    -- successors 2424 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/word_access/word_access_0/rr
      -- 
    split_ack_9413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_gather_scatter_ack_0, ack => cp_elements(2423)); -- 
    rr_9420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2423), ack => ptr_deref_1972_store_0_req_0); -- 
    -- CP-element group 2424 transition  input  no-bypass 
    -- predecessors 2423 
    -- successors 2415 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_request/word_access/word_access_0/ra
      -- 
    ra_9421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_0_ack_0, ack => cp_elements(2424)); -- 
    -- CP-element group 2425 transition  output  bypass 
    -- predecessors 2415 
    -- successors 2426 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2425) <= cp_elements(2415);
    cr_9431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2425), ack => ptr_deref_1972_store_0_req_1); -- 
    -- CP-element group 2426 transition  input  no-bypass 
    -- predecessors 2425 
    -- successors 2416 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1972_complete/word_access/word_access_0/ca
      -- 
    ca_9432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_0_ack_1, ack => cp_elements(2426)); -- 
    -- CP-element group 2427 join  transition  no-bypass 
    -- predecessors 2428 2431 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1978_completed_
      -- 
    cpelement_group_2427 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2428);
      predecessors(1) <= cp_elements(2431);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2427)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2427),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2428 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2427 2429 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1978_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1978_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1977_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1977_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1977_completed_
      -- 
    cp_elements(2428) <= cp_elements(2351);
    -- CP-element group 2429 join  fork  transition  no-bypass 
    -- predecessors 2415 2428 2432 2436 
    -- successors 2430 2437 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_trigger_
      -- 
    cpelement_group_2429 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2415);
      predecessors(1) <= cp_elements(2428);
      predecessors(2) <= cp_elements(2432);
      predecessors(3) <= cp_elements(2436);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2429)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2429),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2430 join  fork  transition  bypass 
    -- predecessors 2429 2439 
    -- successors 2431 2440 2444 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_active_
      -- 
    cpelement_group_2430 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2429);
      predecessors(1) <= cp_elements(2439);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2430)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2430),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2431 join  transition  bypass 
    -- predecessors 2430 2441 
    -- successors 2427 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_completed_
      -- 
    cpelement_group_2431 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2430);
      predecessors(1) <= cp_elements(2441);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2431)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2431),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2432 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2429 2433 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1975_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1975_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1975_completed_
      -- 
    cp_elements(2432) <= cp_elements(2351);
    -- CP-element group 2433 transition  output  bypass 
    -- predecessors 2432 
    -- successors 2434 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_addr_resize/base_resize_req
      -- 
    cp_elements(2433) <= cp_elements(2432);
    base_resize_req_9452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2433), ack => ptr_deref_1976_base_resize_req_0); -- 
    -- CP-element group 2434 transition  input  output  no-bypass 
    -- predecessors 2433 
    -- successors 2435 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_addr_resize/$exit
      -- 
    base_resize_ack_9453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1976_base_resize_ack_0, ack => cp_elements(2434)); -- 
    sum_rename_req_9457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2434), ack => ptr_deref_1976_root_address_inst_req_0); -- 
    -- CP-element group 2435 transition  input  output  no-bypass 
    -- predecessors 2434 
    -- successors 2436 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_word_addrgen/root_register_req
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_base_plus_offset/$exit
      -- 
    sum_rename_ack_9458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1976_root_address_inst_ack_0, ack => cp_elements(2435)); -- 
    root_register_req_9462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2435), ack => ptr_deref_1976_addr_0_req_0); -- 
    -- CP-element group 2436 transition  input  no-bypass 
    -- predecessors 2435 
    -- successors 2429 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_word_addrgen/root_register_ack
      -- 
    root_register_ack_9463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1976_addr_0_ack_0, ack => cp_elements(2436)); -- 
    -- CP-element group 2437 transition  output  bypass 
    -- predecessors 2429 
    -- successors 2438 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/split_req
      -- 
    cp_elements(2437) <= cp_elements(2429);
    split_req_9467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2437), ack => ptr_deref_1976_gather_scatter_req_0); -- 
    -- CP-element group 2438 transition  input  output  no-bypass 
    -- predecessors 2437 
    -- successors 2439 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/split_ack
      -- 
    split_ack_9468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1976_gather_scatter_ack_0, ack => cp_elements(2438)); -- 
    rr_9475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2438), ack => ptr_deref_1976_store_0_req_0); -- 
    -- CP-element group 2439 transition  input  no-bypass 
    -- predecessors 2438 
    -- successors 2430 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_request/$exit
      -- 
    ra_9476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1976_store_0_ack_0, ack => cp_elements(2439)); -- 
    -- CP-element group 2440 transition  output  bypass 
    -- predecessors 2430 
    -- successors 2441 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/word_access/$entry
      -- 
    cp_elements(2440) <= cp_elements(2430);
    cr_9486_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2440), ack => ptr_deref_1976_store_0_req_1); -- 
    -- CP-element group 2441 transition  input  no-bypass 
    -- predecessors 2440 
    -- successors 2431 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1976_complete/word_access/word_access_0/$exit
      -- 
    ca_9487_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1976_store_0_ack_1, ack => cp_elements(2441)); -- 
    -- CP-element group 2442 join  transition  no-bypass 
    -- predecessors 2443 2446 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1982_completed_
      -- 
    cpelement_group_2442 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2443);
      predecessors(1) <= cp_elements(2446);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2442)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2442),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2443 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2442 2444 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1982_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1982_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1981_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1981_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1981_completed_
      -- 
    cp_elements(2443) <= cp_elements(2351);
    -- CP-element group 2444 join  fork  transition  no-bypass 
    -- predecessors 2430 2443 2447 2451 
    -- successors 2445 2452 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_trigger_
      -- 
    cpelement_group_2444 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2430);
      predecessors(1) <= cp_elements(2443);
      predecessors(2) <= cp_elements(2447);
      predecessors(3) <= cp_elements(2451);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2444)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2444),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2445 join  fork  transition  bypass 
    -- predecessors 2444 2454 
    -- successors 2446 2455 2459 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_active_
      -- 
    cpelement_group_2445 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2444);
      predecessors(1) <= cp_elements(2454);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2445)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2445),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2446 join  transition  bypass 
    -- predecessors 2445 2456 
    -- successors 2442 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_completed_
      -- 
    cpelement_group_2446 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2445);
      predecessors(1) <= cp_elements(2456);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2446)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2446),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2447 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2444 2448 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1979_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1979_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1979_completed_
      -- 
    cp_elements(2447) <= cp_elements(2351);
    -- CP-element group 2448 transition  output  bypass 
    -- predecessors 2447 
    -- successors 2449 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_addr_resize/base_resize_req
      -- 
    cp_elements(2448) <= cp_elements(2447);
    base_resize_req_9507_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2448), ack => ptr_deref_1980_base_resize_req_0); -- 
    -- CP-element group 2449 transition  input  output  no-bypass 
    -- predecessors 2448 
    -- successors 2450 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_addr_resize/$exit
      -- 
    base_resize_ack_9508_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1980_base_resize_ack_0, ack => cp_elements(2449)); -- 
    sum_rename_req_9512_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2449), ack => ptr_deref_1980_root_address_inst_req_0); -- 
    -- CP-element group 2450 transition  input  output  no-bypass 
    -- predecessors 2449 
    -- successors 2451 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9513_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1980_root_address_inst_ack_0, ack => cp_elements(2450)); -- 
    root_register_req_9517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2450), ack => ptr_deref_1980_addr_0_req_0); -- 
    -- CP-element group 2451 transition  input  no-bypass 
    -- predecessors 2450 
    -- successors 2444 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_word_addrgen/root_register_ack
      -- 
    root_register_ack_9518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1980_addr_0_ack_0, ack => cp_elements(2451)); -- 
    -- CP-element group 2452 transition  output  bypass 
    -- predecessors 2444 
    -- successors 2453 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/split_req
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/$entry
      -- 
    cp_elements(2452) <= cp_elements(2444);
    split_req_9522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2452), ack => ptr_deref_1980_gather_scatter_req_0); -- 
    -- CP-element group 2453 transition  input  output  no-bypass 
    -- predecessors 2452 
    -- successors 2454 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/word_access/$entry
      -- 
    split_ack_9523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1980_gather_scatter_ack_0, ack => cp_elements(2453)); -- 
    rr_9530_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2453), ack => ptr_deref_1980_store_0_req_0); -- 
    -- CP-element group 2454 transition  input  no-bypass 
    -- predecessors 2453 
    -- successors 2445 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_request/$exit
      -- 
    ra_9531_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1980_store_0_ack_0, ack => cp_elements(2454)); -- 
    -- CP-element group 2455 transition  output  bypass 
    -- predecessors 2445 
    -- successors 2456 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/word_access/$entry
      -- 
    cp_elements(2455) <= cp_elements(2445);
    cr_9541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2455), ack => ptr_deref_1980_store_0_req_1); -- 
    -- CP-element group 2456 transition  input  no-bypass 
    -- predecessors 2455 
    -- successors 2446 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1980_complete/word_access/word_access_0/ca
      -- 
    ca_9542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1980_store_0_ack_1, ack => cp_elements(2456)); -- 
    -- CP-element group 2457 join  transition  no-bypass 
    -- predecessors 2458 2461 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1986_completed_
      -- 
    cpelement_group_2457 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2458);
      predecessors(1) <= cp_elements(2461);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2457)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2457),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2458 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2457 2459 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1985_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1986_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1986_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1985_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1985_completed_
      -- 
    cp_elements(2458) <= cp_elements(2351);
    -- CP-element group 2459 join  fork  transition  no-bypass 
    -- predecessors 2445 2458 2462 2466 
    -- successors 2460 2467 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_trigger_
      -- 
    cpelement_group_2459 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2445);
      predecessors(1) <= cp_elements(2458);
      predecessors(2) <= cp_elements(2462);
      predecessors(3) <= cp_elements(2466);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2459)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2459),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2460 join  fork  transition  bypass 
    -- predecessors 2459 2469 
    -- successors 2461 2470 2474 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_active_
      -- 
    cpelement_group_2460 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2459);
      predecessors(1) <= cp_elements(2469);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2460)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2460),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2461 join  transition  bypass 
    -- predecessors 2460 2471 
    -- successors 2457 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_completed_
      -- 
    cpelement_group_2461 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2460);
      predecessors(1) <= cp_elements(2471);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2461)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2461),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2462 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2459 2463 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1983_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1983_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1983_completed_
      -- 
    cp_elements(2462) <= cp_elements(2351);
    -- CP-element group 2463 transition  output  bypass 
    -- predecessors 2462 
    -- successors 2464 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_addr_resize/base_resize_req
      -- 
    cp_elements(2463) <= cp_elements(2462);
    base_resize_req_9562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2463), ack => ptr_deref_1984_base_resize_req_0); -- 
    -- CP-element group 2464 transition  input  output  no-bypass 
    -- predecessors 2463 
    -- successors 2465 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1984_base_resize_ack_0, ack => cp_elements(2464)); -- 
    sum_rename_req_9567_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2464), ack => ptr_deref_1984_root_address_inst_req_0); -- 
    -- CP-element group 2465 transition  input  output  no-bypass 
    -- predecessors 2464 
    -- successors 2466 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9568_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1984_root_address_inst_ack_0, ack => cp_elements(2465)); -- 
    root_register_req_9572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2465), ack => ptr_deref_1984_addr_0_req_0); -- 
    -- CP-element group 2466 transition  input  no-bypass 
    -- predecessors 2465 
    -- successors 2459 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_word_addrgen/root_register_ack
      -- 
    root_register_ack_9573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1984_addr_0_ack_0, ack => cp_elements(2466)); -- 
    -- CP-element group 2467 transition  output  bypass 
    -- predecessors 2459 
    -- successors 2468 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/split_req
      -- 
    cp_elements(2467) <= cp_elements(2459);
    split_req_9577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2467), ack => ptr_deref_1984_gather_scatter_req_0); -- 
    -- CP-element group 2468 transition  input  output  no-bypass 
    -- predecessors 2467 
    -- successors 2469 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/word_access/word_access_0/rr
      -- 
    split_ack_9578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1984_gather_scatter_ack_0, ack => cp_elements(2468)); -- 
    rr_9585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2468), ack => ptr_deref_1984_store_0_req_0); -- 
    -- CP-element group 2469 transition  input  no-bypass 
    -- predecessors 2468 
    -- successors 2460 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_request/word_access/word_access_0/ra
      -- 
    ra_9586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1984_store_0_ack_0, ack => cp_elements(2469)); -- 
    -- CP-element group 2470 transition  output  bypass 
    -- predecessors 2460 
    -- successors 2471 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2470) <= cp_elements(2460);
    cr_9596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2470), ack => ptr_deref_1984_store_0_req_1); -- 
    -- CP-element group 2471 transition  input  no-bypass 
    -- predecessors 2470 
    -- successors 2461 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1984_complete/word_access/word_access_0/ca
      -- 
    ca_9597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1984_store_0_ack_1, ack => cp_elements(2471)); -- 
    -- CP-element group 2472 join  transition  no-bypass 
    -- predecessors 2473 2476 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1990_completed_
      -- 
    cpelement_group_2472 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2473);
      predecessors(1) <= cp_elements(2476);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2472)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2472),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2473 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2472 2474 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1990_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1990_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1989_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1989_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1989_completed_
      -- 
    cp_elements(2473) <= cp_elements(2351);
    -- CP-element group 2474 join  fork  transition  no-bypass 
    -- predecessors 2460 2473 2477 2481 
    -- successors 2475 2482 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_trigger_
      -- 
    cpelement_group_2474 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2460);
      predecessors(1) <= cp_elements(2473);
      predecessors(2) <= cp_elements(2477);
      predecessors(3) <= cp_elements(2481);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2474)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2474),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2475 join  fork  transition  bypass 
    -- predecessors 2474 2484 
    -- successors 2476 2485 2489 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_active_
      -- 
    cpelement_group_2475 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2474);
      predecessors(1) <= cp_elements(2484);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2475)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2475),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2476 join  transition  bypass 
    -- predecessors 2475 2486 
    -- successors 2472 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_completed_
      -- 
    cpelement_group_2476 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2475);
      predecessors(1) <= cp_elements(2486);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2476)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2476),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2477 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2474 2478 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1987_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1987_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1987_completed_
      -- 
    cp_elements(2477) <= cp_elements(2351);
    -- CP-element group 2478 transition  output  bypass 
    -- predecessors 2477 
    -- successors 2479 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_addr_resize/base_resize_req
      -- 
    cp_elements(2478) <= cp_elements(2477);
    base_resize_req_9617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2478), ack => ptr_deref_1988_base_resize_req_0); -- 
    -- CP-element group 2479 transition  input  output  no-bypass 
    -- predecessors 2478 
    -- successors 2480 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_base_resize_ack_0, ack => cp_elements(2479)); -- 
    sum_rename_req_9622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2479), ack => ptr_deref_1988_root_address_inst_req_0); -- 
    -- CP-element group 2480 transition  input  output  no-bypass 
    -- predecessors 2479 
    -- successors 2481 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_root_address_inst_ack_0, ack => cp_elements(2480)); -- 
    root_register_req_9627_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2480), ack => ptr_deref_1988_addr_0_req_0); -- 
    -- CP-element group 2481 transition  input  no-bypass 
    -- predecessors 2480 
    -- successors 2474 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_word_addrgen/root_register_ack
      -- 
    root_register_ack_9628_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_addr_0_ack_0, ack => cp_elements(2481)); -- 
    -- CP-element group 2482 transition  output  bypass 
    -- predecessors 2474 
    -- successors 2483 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/split_req
      -- 
    cp_elements(2482) <= cp_elements(2474);
    split_req_9632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2482), ack => ptr_deref_1988_gather_scatter_req_0); -- 
    -- CP-element group 2483 transition  input  output  no-bypass 
    -- predecessors 2482 
    -- successors 2484 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/word_access/word_access_0/rr
      -- 
    split_ack_9633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_gather_scatter_ack_0, ack => cp_elements(2483)); -- 
    rr_9640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2483), ack => ptr_deref_1988_store_0_req_0); -- 
    -- CP-element group 2484 transition  input  no-bypass 
    -- predecessors 2483 
    -- successors 2475 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_request/word_access/word_access_0/ra
      -- 
    ra_9641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_store_0_ack_0, ack => cp_elements(2484)); -- 
    -- CP-element group 2485 transition  output  bypass 
    -- predecessors 2475 
    -- successors 2486 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2485) <= cp_elements(2475);
    cr_9651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2485), ack => ptr_deref_1988_store_0_req_1); -- 
    -- CP-element group 2486 transition  input  no-bypass 
    -- predecessors 2485 
    -- successors 2476 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1988_complete/word_access/word_access_0/ca
      -- 
    ca_9652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1988_store_0_ack_1, ack => cp_elements(2486)); -- 
    -- CP-element group 2487 join  transition  no-bypass 
    -- predecessors 2488 2491 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1994_completed_
      -- 
    cpelement_group_2487 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2488);
      predecessors(1) <= cp_elements(2491);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2487)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2487),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2488 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2487 2489 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1994_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1994_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1993_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1993_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1993_completed_
      -- 
    cp_elements(2488) <= cp_elements(2351);
    -- CP-element group 2489 join  fork  transition  no-bypass 
    -- predecessors 2475 2488 2492 2496 
    -- successors 2490 2497 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_trigger_
      -- 
    cpelement_group_2489 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2475);
      predecessors(1) <= cp_elements(2488);
      predecessors(2) <= cp_elements(2492);
      predecessors(3) <= cp_elements(2496);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2489)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2489),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2490 join  fork  transition  bypass 
    -- predecessors 2489 2499 
    -- successors 2491 2500 2504 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_active_
      -- 
    cpelement_group_2490 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2489);
      predecessors(1) <= cp_elements(2499);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2490)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2490),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2491 join  transition  bypass 
    -- predecessors 2490 2501 
    -- successors 2487 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_completed_
      -- 
    cpelement_group_2491 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2490);
      predecessors(1) <= cp_elements(2501);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2491)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2491),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2492 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2489 2493 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1991_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1991_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1991_completed_
      -- 
    cp_elements(2492) <= cp_elements(2351);
    -- CP-element group 2493 transition  output  bypass 
    -- predecessors 2492 
    -- successors 2494 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_addr_resize/base_resize_req
      -- 
    cp_elements(2493) <= cp_elements(2492);
    base_resize_req_9672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2493), ack => ptr_deref_1992_base_resize_req_0); -- 
    -- CP-element group 2494 transition  input  output  no-bypass 
    -- predecessors 2493 
    -- successors 2495 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1992_base_resize_ack_0, ack => cp_elements(2494)); -- 
    sum_rename_req_9677_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2494), ack => ptr_deref_1992_root_address_inst_req_0); -- 
    -- CP-element group 2495 transition  input  output  no-bypass 
    -- predecessors 2494 
    -- successors 2496 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9678_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1992_root_address_inst_ack_0, ack => cp_elements(2495)); -- 
    root_register_req_9682_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2495), ack => ptr_deref_1992_addr_0_req_0); -- 
    -- CP-element group 2496 transition  input  no-bypass 
    -- predecessors 2495 
    -- successors 2489 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_word_addrgen/root_register_ack
      -- 
    root_register_ack_9683_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1992_addr_0_ack_0, ack => cp_elements(2496)); -- 
    -- CP-element group 2497 transition  output  bypass 
    -- predecessors 2489 
    -- successors 2498 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/split_req
      -- 
    cp_elements(2497) <= cp_elements(2489);
    split_req_9687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2497), ack => ptr_deref_1992_gather_scatter_req_0); -- 
    -- CP-element group 2498 transition  input  output  no-bypass 
    -- predecessors 2497 
    -- successors 2499 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/word_access/word_access_0/rr
      -- 
    split_ack_9688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1992_gather_scatter_ack_0, ack => cp_elements(2498)); -- 
    rr_9695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2498), ack => ptr_deref_1992_store_0_req_0); -- 
    -- CP-element group 2499 transition  input  no-bypass 
    -- predecessors 2498 
    -- successors 2490 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_request/word_access/word_access_0/ra
      -- 
    ra_9696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1992_store_0_ack_0, ack => cp_elements(2499)); -- 
    -- CP-element group 2500 transition  output  bypass 
    -- predecessors 2490 
    -- successors 2501 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2500) <= cp_elements(2490);
    cr_9706_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2500), ack => ptr_deref_1992_store_0_req_1); -- 
    -- CP-element group 2501 transition  input  no-bypass 
    -- predecessors 2500 
    -- successors 2491 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1992_complete/word_access/word_access_0/ca
      -- 
    ca_9707_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1992_store_0_ack_1, ack => cp_elements(2501)); -- 
    -- CP-element group 2502 join  transition  no-bypass 
    -- predecessors 2503 2506 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1998_completed_
      -- 
    cpelement_group_2502 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2503);
      predecessors(1) <= cp_elements(2506);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2502)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2502),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2503 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2502 2504 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1998_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_1998_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1997_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1997_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1997_completed_
      -- 
    cp_elements(2503) <= cp_elements(2351);
    -- CP-element group 2504 join  fork  transition  no-bypass 
    -- predecessors 2490 2503 2507 2511 
    -- successors 2505 2512 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_trigger_
      -- 
    cpelement_group_2504 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2490);
      predecessors(1) <= cp_elements(2503);
      predecessors(2) <= cp_elements(2507);
      predecessors(3) <= cp_elements(2511);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2504)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2504),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2505 join  fork  transition  bypass 
    -- predecessors 2504 2514 
    -- successors 2506 2515 2519 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_active_
      -- 
    cpelement_group_2505 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2504);
      predecessors(1) <= cp_elements(2514);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2505)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2505),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2506 join  transition  bypass 
    -- predecessors 2505 2516 
    -- successors 2502 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_completed_
      -- 
    cpelement_group_2506 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2505);
      predecessors(1) <= cp_elements(2516);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2506)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2506),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2507 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2504 2508 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1995_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1995_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1995_completed_
      -- 
    cp_elements(2507) <= cp_elements(2351);
    -- CP-element group 2508 transition  output  bypass 
    -- predecessors 2507 
    -- successors 2509 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_addr_resize/base_resize_req
      -- 
    cp_elements(2508) <= cp_elements(2507);
    base_resize_req_9727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2508), ack => ptr_deref_1996_base_resize_req_0); -- 
    -- CP-element group 2509 transition  input  output  no-bypass 
    -- predecessors 2508 
    -- successors 2510 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9728_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1996_base_resize_ack_0, ack => cp_elements(2509)); -- 
    sum_rename_req_9732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2509), ack => ptr_deref_1996_root_address_inst_req_0); -- 
    -- CP-element group 2510 transition  input  output  no-bypass 
    -- predecessors 2509 
    -- successors 2511 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1996_root_address_inst_ack_0, ack => cp_elements(2510)); -- 
    root_register_req_9737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2510), ack => ptr_deref_1996_addr_0_req_0); -- 
    -- CP-element group 2511 transition  input  no-bypass 
    -- predecessors 2510 
    -- successors 2504 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_word_addrgen/root_register_ack
      -- 
    root_register_ack_9738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1996_addr_0_ack_0, ack => cp_elements(2511)); -- 
    -- CP-element group 2512 transition  output  bypass 
    -- predecessors 2504 
    -- successors 2513 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/split_req
      -- 
    cp_elements(2512) <= cp_elements(2504);
    split_req_9742_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2512), ack => ptr_deref_1996_gather_scatter_req_0); -- 
    -- CP-element group 2513 transition  input  output  no-bypass 
    -- predecessors 2512 
    -- successors 2514 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/word_access/word_access_0/rr
      -- 
    split_ack_9743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1996_gather_scatter_ack_0, ack => cp_elements(2513)); -- 
    rr_9750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2513), ack => ptr_deref_1996_store_0_req_0); -- 
    -- CP-element group 2514 transition  input  no-bypass 
    -- predecessors 2513 
    -- successors 2505 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_request/word_access/word_access_0/ra
      -- 
    ra_9751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1996_store_0_ack_0, ack => cp_elements(2514)); -- 
    -- CP-element group 2515 transition  output  bypass 
    -- predecessors 2505 
    -- successors 2516 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2515) <= cp_elements(2505);
    cr_9761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2515), ack => ptr_deref_1996_store_0_req_1); -- 
    -- CP-element group 2516 transition  input  no-bypass 
    -- predecessors 2515 
    -- successors 2506 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_1996_complete/word_access/word_access_0/ca
      -- 
    ca_9762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1996_store_0_ack_1, ack => cp_elements(2516)); -- 
    -- CP-element group 2517 join  transition  no-bypass 
    -- predecessors 2518 2521 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2002_completed_
      -- 
    cpelement_group_2517 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2518);
      predecessors(1) <= cp_elements(2521);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2517)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2517),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2518 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2517 2519 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2002_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2002_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2001_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2001_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2001_completed_
      -- 
    cp_elements(2518) <= cp_elements(2351);
    -- CP-element group 2519 join  fork  transition  no-bypass 
    -- predecessors 2505 2518 2522 2526 
    -- successors 2520 2527 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_trigger_
      -- 
    cpelement_group_2519 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2505);
      predecessors(1) <= cp_elements(2518);
      predecessors(2) <= cp_elements(2522);
      predecessors(3) <= cp_elements(2526);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2519)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2519),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2520 join  fork  transition  bypass 
    -- predecessors 2519 2529 
    -- successors 2521 2530 2534 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_active_
      -- 
    cpelement_group_2520 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2519);
      predecessors(1) <= cp_elements(2529);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2520)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2520),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2521 join  transition  bypass 
    -- predecessors 2520 2531 
    -- successors 2517 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_completed_
      -- 
    cpelement_group_2521 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2520);
      predecessors(1) <= cp_elements(2531);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2521)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2521),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2522 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2519 2523 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1999_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1999_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_1999_completed_
      -- 
    cp_elements(2522) <= cp_elements(2351);
    -- CP-element group 2523 transition  output  bypass 
    -- predecessors 2522 
    -- successors 2524 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_addr_resize/base_resize_req
      -- 
    cp_elements(2523) <= cp_elements(2522);
    base_resize_req_9782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2523), ack => ptr_deref_2000_base_resize_req_0); -- 
    -- CP-element group 2524 transition  input  output  no-bypass 
    -- predecessors 2523 
    -- successors 2525 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9783_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_base_resize_ack_0, ack => cp_elements(2524)); -- 
    sum_rename_req_9787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2524), ack => ptr_deref_2000_root_address_inst_req_0); -- 
    -- CP-element group 2525 transition  input  output  no-bypass 
    -- predecessors 2524 
    -- successors 2526 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_root_address_inst_ack_0, ack => cp_elements(2525)); -- 
    root_register_req_9792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2525), ack => ptr_deref_2000_addr_0_req_0); -- 
    -- CP-element group 2526 transition  input  no-bypass 
    -- predecessors 2525 
    -- successors 2519 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_word_addrgen/root_register_ack
      -- 
    root_register_ack_9793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_addr_0_ack_0, ack => cp_elements(2526)); -- 
    -- CP-element group 2527 transition  output  bypass 
    -- predecessors 2519 
    -- successors 2528 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/split_req
      -- 
    cp_elements(2527) <= cp_elements(2519);
    split_req_9797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2527), ack => ptr_deref_2000_gather_scatter_req_0); -- 
    -- CP-element group 2528 transition  input  output  no-bypass 
    -- predecessors 2527 
    -- successors 2529 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/word_access/word_access_0/rr
      -- 
    split_ack_9798_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_gather_scatter_ack_0, ack => cp_elements(2528)); -- 
    rr_9805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2528), ack => ptr_deref_2000_store_0_req_0); -- 
    -- CP-element group 2529 transition  input  no-bypass 
    -- predecessors 2528 
    -- successors 2520 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_request/word_access/word_access_0/ra
      -- 
    ra_9806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_store_0_ack_0, ack => cp_elements(2529)); -- 
    -- CP-element group 2530 transition  output  bypass 
    -- predecessors 2520 
    -- successors 2531 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2530) <= cp_elements(2520);
    cr_9816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2530), ack => ptr_deref_2000_store_0_req_1); -- 
    -- CP-element group 2531 transition  input  no-bypass 
    -- predecessors 2530 
    -- successors 2521 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2000_complete/word_access/word_access_0/ca
      -- 
    ca_9817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2000_store_0_ack_1, ack => cp_elements(2531)); -- 
    -- CP-element group 2532 join  transition  no-bypass 
    -- predecessors 2533 2536 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2006_completed_
      -- 
    cpelement_group_2532 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2533);
      predecessors(1) <= cp_elements(2536);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2532)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2532),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2533 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2532 2534 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2005_completed_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2006_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2006_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2005_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2005_active_
      -- 
    cp_elements(2533) <= cp_elements(2351);
    -- CP-element group 2534 join  fork  transition  no-bypass 
    -- predecessors 2520 2533 2537 2541 
    -- successors 2535 2542 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_trigger_
      -- 
    cpelement_group_2534 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2520);
      predecessors(1) <= cp_elements(2533);
      predecessors(2) <= cp_elements(2537);
      predecessors(3) <= cp_elements(2541);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2534)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2534),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2535 join  fork  transition  bypass 
    -- predecessors 2534 2544 
    -- successors 2536 2545 2549 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_active_
      -- 
    cpelement_group_2535 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2534);
      predecessors(1) <= cp_elements(2544);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2535)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2535),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2536 join  transition  bypass 
    -- predecessors 2535 2546 
    -- successors 2532 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_completed_
      -- 
    cpelement_group_2536 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2535);
      predecessors(1) <= cp_elements(2546);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2536)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2536),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2537 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2534 2538 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2003_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2003_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2003_completed_
      -- 
    cp_elements(2537) <= cp_elements(2351);
    -- CP-element group 2538 transition  output  bypass 
    -- predecessors 2537 
    -- successors 2539 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_addr_resize/base_resize_req
      -- 
    cp_elements(2538) <= cp_elements(2537);
    base_resize_req_9837_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2538), ack => ptr_deref_2004_base_resize_req_0); -- 
    -- CP-element group 2539 transition  input  output  no-bypass 
    -- predecessors 2538 
    -- successors 2540 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9838_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2004_base_resize_ack_0, ack => cp_elements(2539)); -- 
    sum_rename_req_9842_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2539), ack => ptr_deref_2004_root_address_inst_req_0); -- 
    -- CP-element group 2540 transition  input  output  no-bypass 
    -- predecessors 2539 
    -- successors 2541 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9843_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2004_root_address_inst_ack_0, ack => cp_elements(2540)); -- 
    root_register_req_9847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2540), ack => ptr_deref_2004_addr_0_req_0); -- 
    -- CP-element group 2541 transition  input  no-bypass 
    -- predecessors 2540 
    -- successors 2534 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_word_addrgen/root_register_ack
      -- 
    root_register_ack_9848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2004_addr_0_ack_0, ack => cp_elements(2541)); -- 
    -- CP-element group 2542 transition  output  bypass 
    -- predecessors 2534 
    -- successors 2543 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/split_req
      -- 
    cp_elements(2542) <= cp_elements(2534);
    split_req_9852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2542), ack => ptr_deref_2004_gather_scatter_req_0); -- 
    -- CP-element group 2543 transition  input  output  no-bypass 
    -- predecessors 2542 
    -- successors 2544 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/word_access/word_access_0/rr
      -- 
    split_ack_9853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2004_gather_scatter_ack_0, ack => cp_elements(2543)); -- 
    rr_9860_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2543), ack => ptr_deref_2004_store_0_req_0); -- 
    -- CP-element group 2544 transition  input  no-bypass 
    -- predecessors 2543 
    -- successors 2535 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_request/word_access/word_access_0/ra
      -- 
    ra_9861_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2004_store_0_ack_0, ack => cp_elements(2544)); -- 
    -- CP-element group 2545 transition  output  bypass 
    -- predecessors 2535 
    -- successors 2546 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2545) <= cp_elements(2535);
    cr_9871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2545), ack => ptr_deref_2004_store_0_req_1); -- 
    -- CP-element group 2546 transition  input  no-bypass 
    -- predecessors 2545 
    -- successors 2536 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2004_complete/word_access/word_access_0/ca
      -- 
    ca_9872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2004_store_0_ack_1, ack => cp_elements(2546)); -- 
    -- CP-element group 2547 join  transition  no-bypass 
    -- predecessors 2548 2551 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2010_completed_
      -- 
    cpelement_group_2547 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2548);
      predecessors(1) <= cp_elements(2551);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2547)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2547),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2548 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2547 2549 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2010_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2010_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2009_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2009_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2009_completed_
      -- 
    cp_elements(2548) <= cp_elements(2351);
    -- CP-element group 2549 join  fork  transition  no-bypass 
    -- predecessors 2535 2548 2552 2556 
    -- successors 2550 2557 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_trigger_
      -- 
    cpelement_group_2549 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2535);
      predecessors(1) <= cp_elements(2548);
      predecessors(2) <= cp_elements(2552);
      predecessors(3) <= cp_elements(2556);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2549)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2549),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2550 join  fork  transition  bypass 
    -- predecessors 2549 2559 
    -- successors 2551 2560 2564 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_active_
      -- 
    cpelement_group_2550 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2549);
      predecessors(1) <= cp_elements(2559);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2550)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2550),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2551 join  transition  bypass 
    -- predecessors 2550 2561 
    -- successors 2547 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_completed_
      -- 
    cpelement_group_2551 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2550);
      predecessors(1) <= cp_elements(2561);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2551)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2551),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2552 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2549 2553 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2007_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2007_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2007_completed_
      -- 
    cp_elements(2552) <= cp_elements(2351);
    -- CP-element group 2553 transition  output  bypass 
    -- predecessors 2552 
    -- successors 2554 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_addr_resize/base_resize_req
      -- 
    cp_elements(2553) <= cp_elements(2552);
    base_resize_req_9892_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2553), ack => ptr_deref_2008_base_resize_req_0); -- 
    -- CP-element group 2554 transition  input  output  no-bypass 
    -- predecessors 2553 
    -- successors 2555 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9893_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2008_base_resize_ack_0, ack => cp_elements(2554)); -- 
    sum_rename_req_9897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2554), ack => ptr_deref_2008_root_address_inst_req_0); -- 
    -- CP-element group 2555 transition  input  output  no-bypass 
    -- predecessors 2554 
    -- successors 2556 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2008_root_address_inst_ack_0, ack => cp_elements(2555)); -- 
    root_register_req_9902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2555), ack => ptr_deref_2008_addr_0_req_0); -- 
    -- CP-element group 2556 transition  input  no-bypass 
    -- predecessors 2555 
    -- successors 2549 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_word_addrgen/root_register_ack
      -- 
    root_register_ack_9903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2008_addr_0_ack_0, ack => cp_elements(2556)); -- 
    -- CP-element group 2557 transition  output  bypass 
    -- predecessors 2549 
    -- successors 2558 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/split_req
      -- 
    cp_elements(2557) <= cp_elements(2549);
    split_req_9907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2557), ack => ptr_deref_2008_gather_scatter_req_0); -- 
    -- CP-element group 2558 transition  input  output  no-bypass 
    -- predecessors 2557 
    -- successors 2559 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/word_access/word_access_0/rr
      -- 
    split_ack_9908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2008_gather_scatter_ack_0, ack => cp_elements(2558)); -- 
    rr_9915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2558), ack => ptr_deref_2008_store_0_req_0); -- 
    -- CP-element group 2559 transition  input  no-bypass 
    -- predecessors 2558 
    -- successors 2550 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_request/word_access/word_access_0/ra
      -- 
    ra_9916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2008_store_0_ack_0, ack => cp_elements(2559)); -- 
    -- CP-element group 2560 transition  output  bypass 
    -- predecessors 2550 
    -- successors 2561 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2560) <= cp_elements(2550);
    cr_9926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2560), ack => ptr_deref_2008_store_0_req_1); -- 
    -- CP-element group 2561 transition  input  no-bypass 
    -- predecessors 2560 
    -- successors 2551 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2008_complete/word_access/word_access_0/ca
      -- 
    ca_9927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2008_store_0_ack_1, ack => cp_elements(2561)); -- 
    -- CP-element group 2562 join  transition  no-bypass 
    -- predecessors 2563 2566 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2014_completed_
      -- 
    cpelement_group_2562 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2563);
      predecessors(1) <= cp_elements(2566);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2562)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2562),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2563 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2562 2564 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2014_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2014_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2013_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2013_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2013_completed_
      -- 
    cp_elements(2563) <= cp_elements(2351);
    -- CP-element group 2564 join  fork  transition  no-bypass 
    -- predecessors 2550 2563 2567 2571 
    -- successors 2565 2572 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_trigger_
      -- 
    cpelement_group_2564 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2550);
      predecessors(1) <= cp_elements(2563);
      predecessors(2) <= cp_elements(2567);
      predecessors(3) <= cp_elements(2571);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2564)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2564),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2565 join  fork  transition  bypass 
    -- predecessors 2564 2574 
    -- successors 2566 2575 2579 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_active_
      -- 
    cpelement_group_2565 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2564);
      predecessors(1) <= cp_elements(2574);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2565)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2565),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2566 join  transition  bypass 
    -- predecessors 2565 2576 
    -- successors 2562 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_completed_
      -- 
    cpelement_group_2566 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2565);
      predecessors(1) <= cp_elements(2576);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2566)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2566),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2567 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2564 2568 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2011_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2011_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2011_completed_
      -- 
    cp_elements(2567) <= cp_elements(2351);
    -- CP-element group 2568 transition  output  bypass 
    -- predecessors 2567 
    -- successors 2569 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_addr_resize/base_resize_req
      -- 
    cp_elements(2568) <= cp_elements(2567);
    base_resize_req_9947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2568), ack => ptr_deref_2012_base_resize_req_0); -- 
    -- CP-element group 2569 transition  input  output  no-bypass 
    -- predecessors 2568 
    -- successors 2570 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_9948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2012_base_resize_ack_0, ack => cp_elements(2569)); -- 
    sum_rename_req_9952_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2569), ack => ptr_deref_2012_root_address_inst_req_0); -- 
    -- CP-element group 2570 transition  input  output  no-bypass 
    -- predecessors 2569 
    -- successors 2571 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_word_addrgen/root_register_req
      -- 
    sum_rename_ack_9953_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2012_root_address_inst_ack_0, ack => cp_elements(2570)); -- 
    root_register_req_9957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2570), ack => ptr_deref_2012_addr_0_req_0); -- 
    -- CP-element group 2571 transition  input  no-bypass 
    -- predecessors 2570 
    -- successors 2564 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_word_addrgen/root_register_ack
      -- 
    root_register_ack_9958_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2012_addr_0_ack_0, ack => cp_elements(2571)); -- 
    -- CP-element group 2572 transition  output  bypass 
    -- predecessors 2564 
    -- successors 2573 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/split_req
      -- 
    cp_elements(2572) <= cp_elements(2564);
    split_req_9962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2572), ack => ptr_deref_2012_gather_scatter_req_0); -- 
    -- CP-element group 2573 transition  input  output  no-bypass 
    -- predecessors 2572 
    -- successors 2574 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/word_access/word_access_0/rr
      -- 
    split_ack_9963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2012_gather_scatter_ack_0, ack => cp_elements(2573)); -- 
    rr_9970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2573), ack => ptr_deref_2012_store_0_req_0); -- 
    -- CP-element group 2574 transition  input  no-bypass 
    -- predecessors 2573 
    -- successors 2565 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_request/word_access/word_access_0/ra
      -- 
    ra_9971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2012_store_0_ack_0, ack => cp_elements(2574)); -- 
    -- CP-element group 2575 transition  output  bypass 
    -- predecessors 2565 
    -- successors 2576 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2575) <= cp_elements(2565);
    cr_9981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2575), ack => ptr_deref_2012_store_0_req_1); -- 
    -- CP-element group 2576 transition  input  no-bypass 
    -- predecessors 2575 
    -- successors 2566 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2012_complete/word_access/word_access_0/ca
      -- 
    ca_9982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2012_store_0_ack_1, ack => cp_elements(2576)); -- 
    -- CP-element group 2577 join  transition  no-bypass 
    -- predecessors 2578 2581 
    -- successors 2605 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2018_completed_
      -- 
    cpelement_group_2577 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2578);
      predecessors(1) <= cp_elements(2581);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2577)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2577),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2578 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2577 2579 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2018_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2018_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2017_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2017_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2017_completed_
      -- 
    cp_elements(2578) <= cp_elements(2351);
    -- CP-element group 2579 join  fork  transition  no-bypass 
    -- predecessors 2565 2578 2582 2586 
    -- successors 2580 2587 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_trigger_
      -- 
    cpelement_group_2579 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2565);
      predecessors(1) <= cp_elements(2578);
      predecessors(2) <= cp_elements(2582);
      predecessors(3) <= cp_elements(2586);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2579)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2579),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2580 join  fork  transition  bypass 
    -- predecessors 2579 2589 
    -- successors 2581 2590 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_active_
      -- 
    cpelement_group_2580 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2579);
      predecessors(1) <= cp_elements(2589);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2580)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2580),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2581 join  transition  bypass 
    -- predecessors 2580 2591 
    -- successors 2577 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_completed_
      -- 
    cpelement_group_2581 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2580);
      predecessors(1) <= cp_elements(2591);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2581)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2581),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2582 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2579 2583 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2015_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2015_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2015_completed_
      -- 
    cp_elements(2582) <= cp_elements(2351);
    -- CP-element group 2583 transition  output  bypass 
    -- predecessors 2582 
    -- successors 2584 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_addr_resize/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_addr_resize/base_resize_req
      -- 
    cp_elements(2583) <= cp_elements(2582);
    base_resize_req_10002_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2583), ack => ptr_deref_2016_base_resize_req_0); -- 
    -- CP-element group 2584 transition  input  output  no-bypass 
    -- predecessors 2583 
    -- successors 2585 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_address_resized
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_addr_resize/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_plus_offset/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_10003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2016_base_resize_ack_0, ack => cp_elements(2584)); -- 
    sum_rename_req_10007_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2584), ack => ptr_deref_2016_root_address_inst_req_0); -- 
    -- CP-element group 2585 transition  input  output  no-bypass 
    -- predecessors 2584 
    -- successors 2586 
    -- members (5) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_root_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_plus_offset/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_word_addrgen/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_word_addrgen/root_register_req
      -- 
    sum_rename_ack_10008_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2016_root_address_inst_ack_0, ack => cp_elements(2585)); -- 
    root_register_req_10012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2585), ack => ptr_deref_2016_addr_0_req_0); -- 
    -- CP-element group 2586 transition  input  no-bypass 
    -- predecessors 2585 
    -- successors 2579 
    -- members (3) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_word_address_calculated
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_word_addrgen/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_word_addrgen/root_register_ack
      -- 
    root_register_ack_10013_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2016_addr_0_ack_0, ack => cp_elements(2586)); -- 
    -- CP-element group 2587 transition  output  bypass 
    -- predecessors 2579 
    -- successors 2588 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/split_req
      -- 
    cp_elements(2587) <= cp_elements(2579);
    split_req_10017_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2587), ack => ptr_deref_2016_gather_scatter_req_0); -- 
    -- CP-element group 2588 transition  input  output  no-bypass 
    -- predecessors 2587 
    -- successors 2589 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/split_ack
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/word_access/word_access_0/rr
      -- 
    split_ack_10018_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2016_gather_scatter_ack_0, ack => cp_elements(2588)); -- 
    rr_10025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2588), ack => ptr_deref_2016_store_0_req_0); -- 
    -- CP-element group 2589 transition  input  no-bypass 
    -- predecessors 2588 
    -- successors 2580 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_request/word_access/word_access_0/ra
      -- 
    ra_10026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2016_store_0_ack_0, ack => cp_elements(2589)); -- 
    -- CP-element group 2590 transition  output  bypass 
    -- predecessors 2580 
    -- successors 2591 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/word_access/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/word_access/word_access_0/cr
      -- 
    cp_elements(2590) <= cp_elements(2580);
    cr_10036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2590), ack => ptr_deref_2016_store_0_req_1); -- 
    -- CP-element group 2591 transition  input  no-bypass 
    -- predecessors 2590 
    -- successors 2581 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/word_access/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/ptr_deref_2016_complete/word_access/word_access_0/ca
      -- 
    ca_10037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2016_store_0_ack_1, ack => cp_elements(2591)); -- 
    -- CP-element group 2592 join  fork  transition  no-bypass 
    -- predecessors 2594 2596 
    -- successors 2593 2597 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_active_
      -- 
    cpelement_group_2592 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2594);
      predecessors(1) <= cp_elements(2596);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2592)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2592),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2593 join  fork  transition  bypass 
    -- predecessors 2592 2598 
    -- successors 2599 2601 
    -- members (8) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2024_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2024_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2024_completed_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_completed_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2026_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2026_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2026_completed_
      -- 
    cpelement_group_2593 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2592);
      predecessors(1) <= cp_elements(2598);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2593)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2593),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2594 fork  transition  bypass 
    -- predecessors 2351 
    -- successors 2592 2595 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2020_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2020_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/simple_obj_ref_2020_completed_
      -- 
    cp_elements(2594) <= cp_elements(2351);
    -- CP-element group 2595 transition  output  bypass 
    -- predecessors 2594 
    -- successors 2596 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Sample/rr
      -- 
    cp_elements(2595) <= cp_elements(2594);
    rr_10050_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2595), ack => binary_2023_inst_req_0); -- 
    -- CP-element group 2596 transition  input  no-bypass 
    -- predecessors 2595 
    -- successors 2592 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Sample/ra
      -- 
    ra_10051_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2023_inst_ack_0, ack => cp_elements(2596)); -- 
    -- CP-element group 2597 transition  output  bypass 
    -- predecessors 2592 
    -- successors 2598 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Update/cr
      -- 
    cp_elements(2597) <= cp_elements(2592);
    cr_10055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2597), ack => binary_2023_inst_req_1); -- 
    -- CP-element group 2598 transition  input  no-bypass 
    -- predecessors 2597 
    -- successors 2593 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2023_complete_Update/ca
      -- 
    ca_10056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2023_inst_ack_1, ack => cp_elements(2598)); -- 
    -- CP-element group 2599 join  fork  transition  bypass 
    -- predecessors 2593 2602 
    -- successors 2600 2603 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_active_
      -- 
    cpelement_group_2599 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2593);
      predecessors(1) <= cp_elements(2602);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2599)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2599),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2600 join  transition  no-bypass 
    -- predecessors 2599 2604 
    -- successors 2605 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2030_trigger_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2030_active_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/assign_stmt_2030_completed_
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_completed_
      -- 
    cpelement_group_2600 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2599);
      predecessors(1) <= cp_elements(2604);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2600)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2600),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2601 transition  output  bypass 
    -- predecessors 2593 
    -- successors 2602 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Sample/rr
      -- 
    cp_elements(2601) <= cp_elements(2593);
    rr_10069_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2601), ack => binary_2029_inst_req_0); -- 
    -- CP-element group 2602 transition  input  no-bypass 
    -- predecessors 2601 
    -- successors 2599 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Sample/ra
      -- 
    ra_10070_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2029_inst_ack_0, ack => cp_elements(2602)); -- 
    -- CP-element group 2603 transition  output  bypass 
    -- predecessors 2599 
    -- successors 2604 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Update/cr
      -- 
    cp_elements(2603) <= cp_elements(2599);
    cr_10074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2603), ack => binary_2029_inst_req_1); -- 
    -- CP-element group 2604 transition  input  no-bypass 
    -- predecessors 2603 
    -- successors 2600 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/binary_2029_complete_Update/ca
      -- 
    ca_10075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2029_inst_ack_1, ack => cp_elements(2604)); -- 
    -- CP-element group 2605 join  transition  no-bypass 
    -- predecessors 2352 2367 2382 2397 2412 2427 2442 2457 2472 2487 2502 2517 2532 2547 2562 2577 2600 
    -- successors 6 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_1958_to_assign_stmt_2030/$exit
      -- 
    cpelement_group_2605 : Block -- 
      signal predecessors: BooleanArray(16 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2352);
      predecessors(1) <= cp_elements(2367);
      predecessors(2) <= cp_elements(2382);
      predecessors(3) <= cp_elements(2397);
      predecessors(4) <= cp_elements(2412);
      predecessors(5) <= cp_elements(2427);
      predecessors(6) <= cp_elements(2442);
      predecessors(7) <= cp_elements(2457);
      predecessors(8) <= cp_elements(2472);
      predecessors(9) <= cp_elements(2487);
      predecessors(10) <= cp_elements(2502);
      predecessors(11) <= cp_elements(2517);
      predecessors(12) <= cp_elements(2532);
      predecessors(13) <= cp_elements(2547);
      predecessors(14) <= cp_elements(2562);
      predecessors(15) <= cp_elements(2577);
      predecessors(16) <= cp_elements(2600);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2605)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2605),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2606 transition  bypass 
    -- predecessors 6 
    -- successors 2607 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2031_dead_link/$entry
      -- 
    cp_elements(2606) <= cp_elements(6);
    -- CP-element group 2607 transition  dead  bypass 
    -- predecessors 2606 
    -- successors 2608 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2031_dead_link/dead_transition
      -- 
    cp_elements(2607) <= false;
    -- CP-element group 2608 transition  place  bypass 
    -- predecessors 2607 
    -- successors 2774 
    -- members (4) 
      -- 	branch_block_stmt_552/merge_stmt_2037__entry__
      -- 	branch_block_stmt_552/if_stmt_2031__exit__
      -- 	branch_block_stmt_552/if_stmt_2031_dead_link/$exit
      -- 	branch_block_stmt_552/merge_stmt_2037_dead_link/$entry
      -- 
    cp_elements(2608) <= cp_elements(2607);
    -- CP-element group 2609 transition  output  bypass 
    -- predecessors 6 
    -- successors 2610 
    -- members (3) 
      -- 	branch_block_stmt_552/if_stmt_2031_eval_test/$entry
      -- 	branch_block_stmt_552/if_stmt_2031_eval_test/$exit
      -- 	branch_block_stmt_552/if_stmt_2031_eval_test/branch_req
      -- 
    cp_elements(2609) <= cp_elements(6);
    branch_req_10083_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2609), ack => if_stmt_2031_branch_req_0); -- 
    -- CP-element group 2610 branch  place  bypass 
    -- predecessors 2609 
    -- successors 2611 2613 
    -- members (1) 
      -- 	branch_block_stmt_552/simple_obj_ref_2032_place
      -- 
    cp_elements(2610) <= cp_elements(2609);
    -- CP-element group 2611 transition  bypass 
    -- predecessors 2610 
    -- successors 2612 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2031_if_link/$entry
      -- 
    cp_elements(2611) <= cp_elements(2610);
    -- CP-element group 2612 transition  place  input  no-bypass 
    -- predecessors 2611 
    -- successors 7 
    -- members (9) 
      -- 	branch_block_stmt_552/merge_stmt_2037_PhiReqMerge
      -- 	branch_block_stmt_552/if_stmt_2031_if_link/$exit
      -- 	branch_block_stmt_552/if_stmt_2031_if_link/if_choice_transition
      -- 	branch_block_stmt_552/xx_x_crit_edge_xx_x_crit_edge37
      -- 	branch_block_stmt_552/xx_x_crit_edge_xx_x_crit_edge37_PhiReq/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge_xx_x_crit_edge37_PhiReq/$exit
      -- 	branch_block_stmt_552/merge_stmt_2037_PhiAck/$entry
      -- 	branch_block_stmt_552/merge_stmt_2037_PhiAck/$exit
      -- 	branch_block_stmt_552/merge_stmt_2037_PhiAck/dummy
      -- 
    if_choice_transition_10088_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2031_branch_ack_1, ack => cp_elements(2612)); -- 
    -- CP-element group 2613 transition  bypass 
    -- predecessors 2610 
    -- successors 2614 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2031_else_link/$entry
      -- 
    cp_elements(2613) <= cp_elements(2610);
    -- CP-element group 2614 transition  place  input  output  no-bypass 
    -- predecessors 2613 
    -- successors 2640 
    -- members (8) 
      -- 	branch_block_stmt_552/if_stmt_2031_else_link/$exit
      -- 	branch_block_stmt_552/if_stmt_2031_else_link/else_choice_transition
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/req
      -- 
    else_choice_transition_10092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2031_branch_ack_0, ack => cp_elements(2614)); -- 
    req_10217_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2614), ack => type_cast_595_inst_req_0); -- 
    -- CP-element group 2615 join  fork  transition  bypass 
    -- predecessors 7 2618 
    -- successors 2616 2619 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_active_
      -- 
    cpelement_group_2615 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(7);
      predecessors(1) <= cp_elements(2618);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2615)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2615),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2616 join  fork  transition  bypass 
    -- predecessors 2615 2620 
    -- successors 2621 2623 
    -- members (8) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/assign_stmt_2043_trigger_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/assign_stmt_2043_active_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/assign_stmt_2043_completed_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_completed_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_trigger_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/simple_obj_ref_2045_trigger_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/simple_obj_ref_2045_active_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/simple_obj_ref_2045_completed_
      -- 
    cpelement_group_2616 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2615);
      predecessors(1) <= cp_elements(2620);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2616)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2616),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2617 transition  output  bypass 
    -- predecessors 7 
    -- successors 2618 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Sample/rr
      -- 
    cp_elements(2617) <= cp_elements(7);
    rr_10110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2617), ack => binary_2042_inst_req_0); -- 
    -- CP-element group 2618 transition  input  no-bypass 
    -- predecessors 2617 
    -- successors 2615 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Sample/ra
      -- 
    ra_10111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2042_inst_ack_0, ack => cp_elements(2618)); -- 
    -- CP-element group 2619 transition  output  bypass 
    -- predecessors 2615 
    -- successors 2620 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Update/cr
      -- 
    cp_elements(2619) <= cp_elements(2615);
    cr_10115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2619), ack => binary_2042_inst_req_1); -- 
    -- CP-element group 2620 transition  input  no-bypass 
    -- predecessors 2619 
    -- successors 2616 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2042_complete_Update/ca
      -- 
    ca_10116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2042_inst_ack_1, ack => cp_elements(2620)); -- 
    -- CP-element group 2621 join  fork  transition  no-bypass 
    -- predecessors 2616 2624 
    -- successors 2622 2625 
    -- members (1) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_active_
      -- 
    cpelement_group_2621 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2616);
      predecessors(1) <= cp_elements(2624);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2621)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2621),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2622 branch  join  transition  place  no-bypass 
    -- predecessors 2621 2626 
    -- successors 2627 2630 
    -- members (7) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049__exit__
      -- 	branch_block_stmt_552/if_stmt_2050__entry__
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/$exit
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/assign_stmt_2049_trigger_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/assign_stmt_2049_active_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/assign_stmt_2049_completed_
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_completed_
      -- 
    cpelement_group_2622 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2621);
      predecessors(1) <= cp_elements(2626);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2622)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2622),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2623 transition  output  bypass 
    -- predecessors 2616 
    -- successors 2624 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Sample/$entry
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Sample/rr
      -- 
    cp_elements(2623) <= cp_elements(2616);
    rr_10129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2623), ack => binary_2048_inst_req_0); -- 
    -- CP-element group 2624 transition  input  no-bypass 
    -- predecessors 2623 
    -- successors 2621 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Sample/$exit
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Sample/ra
      -- 
    ra_10130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2048_inst_ack_0, ack => cp_elements(2624)); -- 
    -- CP-element group 2625 transition  output  bypass 
    -- predecessors 2621 
    -- successors 2626 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Update/$entry
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Update/cr
      -- 
    cp_elements(2625) <= cp_elements(2621);
    cr_10134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2625), ack => binary_2048_inst_req_1); -- 
    -- CP-element group 2626 transition  input  no-bypass 
    -- predecessors 2625 
    -- successors 2622 
    -- members (2) 
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Update/$exit
      -- 	branch_block_stmt_552/assign_stmt_2043_to_assign_stmt_2049/binary_2048_complete_Update/ca
      -- 
    ca_10135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2048_inst_ack_1, ack => cp_elements(2626)); -- 
    -- CP-element group 2627 transition  bypass 
    -- predecessors 2622 
    -- successors 2628 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2050_dead_link/$entry
      -- 
    cp_elements(2627) <= cp_elements(2622);
    -- CP-element group 2628 transition  dead  bypass 
    -- predecessors 2627 
    -- successors 2629 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2050_dead_link/dead_transition
      -- 
    cp_elements(2628) <= false;
    -- CP-element group 2629 transition  place  bypass 
    -- predecessors 2628 
    -- successors 2776 
    -- members (4) 
      -- 	branch_block_stmt_552/if_stmt_2050__exit__
      -- 	branch_block_stmt_552/merge_stmt_2056__entry__
      -- 	branch_block_stmt_552/if_stmt_2050_dead_link/$exit
      -- 	branch_block_stmt_552/merge_stmt_2056_dead_link/$entry
      -- 
    cp_elements(2629) <= cp_elements(2628);
    -- CP-element group 2630 transition  output  bypass 
    -- predecessors 2622 
    -- successors 2631 
    -- members (3) 
      -- 	branch_block_stmt_552/if_stmt_2050_eval_test/$entry
      -- 	branch_block_stmt_552/if_stmt_2050_eval_test/$exit
      -- 	branch_block_stmt_552/if_stmt_2050_eval_test/branch_req
      -- 
    cp_elements(2630) <= cp_elements(2622);
    branch_req_10143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2630), ack => if_stmt_2050_branch_req_0); -- 
    -- CP-element group 2631 branch  place  bypass 
    -- predecessors 2630 
    -- successors 2632 2634 
    -- members (1) 
      -- 	branch_block_stmt_552/simple_obj_ref_2051_place
      -- 
    cp_elements(2631) <= cp_elements(2630);
    -- CP-element group 2632 transition  bypass 
    -- predecessors 2631 
    -- successors 2633 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2050_if_link/$entry
      -- 
    cp_elements(2632) <= cp_elements(2631);
    -- CP-element group 2633 transition  place  input  no-bypass 
    -- predecessors 2632 
    -- successors 8 
    -- members (9) 
      -- 	branch_block_stmt_552/merge_stmt_2056_PhiReqMerge
      -- 	branch_block_stmt_552/if_stmt_2050_if_link/$exit
      -- 	branch_block_stmt_552/if_stmt_2050_if_link/if_choice_transition
      -- 	branch_block_stmt_552/xx_x_crit_edge37_xx_x_crit_edge40
      -- 	branch_block_stmt_552/xx_x_crit_edge37_xx_x_crit_edge40_PhiReq/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge37_xx_x_crit_edge40_PhiReq/$exit
      -- 	branch_block_stmt_552/merge_stmt_2056_PhiAck/$entry
      -- 	branch_block_stmt_552/merge_stmt_2056_PhiAck/$exit
      -- 	branch_block_stmt_552/merge_stmt_2056_PhiAck/dummy
      -- 
    if_choice_transition_10148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2050_branch_ack_1, ack => cp_elements(2633)); -- 
    -- CP-element group 2634 transition  bypass 
    -- predecessors 2631 
    -- successors 2635 
    -- members (1) 
      -- 	branch_block_stmt_552/if_stmt_2050_else_link/$entry
      -- 
    cp_elements(2634) <= cp_elements(2631);
    -- CP-element group 2635 transition  place  input  output  no-bypass 
    -- predecessors 2634 
    -- successors 2636 
    -- members (8) 
      -- 	branch_block_stmt_552/if_stmt_2050_else_link/$exit
      -- 	branch_block_stmt_552/if_stmt_2050_else_link/else_choice_transition
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/$entry
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/req
      -- 
    else_choice_transition_10152_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2050_branch_ack_0, ack => cp_elements(2635)); -- 
    req_10182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2635), ack => type_cast_561_inst_req_0); -- 
    -- CP-element group 2636 transition  input  output  no-bypass 
    -- predecessors 2635 
    -- successors 2637 
    -- members (6) 
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/ack
      -- 	branch_block_stmt_552/xx_x_crit_edge37_bbx_xnph36_PhiReq/phi_stmt_555/phi_stmt_555_req
      -- 
    ack_10183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => cp_elements(2636)); -- 
    phi_stmt_555_req_10184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2636), ack => phi_stmt_555_req_1); -- 
    -- CP-element group 2637 merge  place  bypass 
    -- predecessors 0 2636 
    -- successors 2638 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_554_PhiReqMerge
      -- 
    cp_elements(2637) <= OrReduce(cp_elements(0) & cp_elements(2636));
    -- CP-element group 2638 transition  bypass 
    -- predecessors 2637 
    -- successors 2639 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_554_PhiAck/$entry
      -- 
    cp_elements(2638) <= cp_elements(2637);
    -- CP-element group 2639 fork  transition  place  input  no-bypass 
    -- predecessors 2638 
    -- successors 9 11 
    -- members (9) 
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_564_completed_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_564_active_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/simple_obj_ref_564_trigger_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586__entry__
      -- 	branch_block_stmt_552/merge_stmt_554__exit__
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/binary_567_trigger_
      -- 	branch_block_stmt_552/assign_stmt_568_to_assign_stmt_586/$entry
      -- 	branch_block_stmt_552/merge_stmt_554_PhiAck/$exit
      -- 	branch_block_stmt_552/merge_stmt_554_PhiAck/phi_stmt_555_ack
      -- 
    phi_stmt_555_ack_10189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_555_ack_0, ack => cp_elements(2639)); -- 
    -- CP-element group 2640 transition  input  output  no-bypass 
    -- predecessors 2614 
    -- successors 2641 
    -- members (6) 
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/$exit
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_sources/type_cast_595/ack
      -- 	branch_block_stmt_552/xx_x_crit_edge_bbx_xnph_PhiReq/phi_stmt_589/phi_stmt_589_req
      -- 
    ack_10218_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_595_inst_ack_0, ack => cp_elements(2640)); -- 
    phi_stmt_589_req_10219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2640), ack => phi_stmt_589_req_1); -- 
    -- CP-element group 2641 merge  place  bypass 
    -- predecessors 1 2640 
    -- successors 2642 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_588_PhiReqMerge
      -- 
    cp_elements(2641) <= OrReduce(cp_elements(1) & cp_elements(2640));
    -- CP-element group 2642 transition  bypass 
    -- predecessors 2641 
    -- successors 2643 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_588_PhiAck/$entry
      -- 
    cp_elements(2642) <= cp_elements(2641);
    -- CP-element group 2643 transition  place  input  no-bypass 
    -- predecessors 2642 
    -- successors 37 
    -- members (4) 
      -- 	branch_block_stmt_552/assign_stmt_602_to_assign_stmt_740__entry__
      -- 	branch_block_stmt_552/merge_stmt_588__exit__
      -- 	branch_block_stmt_552/merge_stmt_588_PhiAck/phi_stmt_589_ack
      -- 	branch_block_stmt_552/merge_stmt_588_PhiAck/$exit
      -- 
    phi_stmt_589_ack_10224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_589_ack_0, ack => cp_elements(2643)); -- 
    -- CP-element group 2644 fork  transition  bypass 
    -- predecessors 2350 
    -- successors 2645 2647 2649 2651 2653 2655 2657 2659 2661 2663 2665 2667 2669 2671 2673 2675 2677 
    -- members (1) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/$entry
      -- 
    cp_elements(2644) <= cp_elements(2350);
    -- CP-element group 2645 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2646 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/$entry
      -- 
    cp_elements(2645) <= cp_elements(2644);
    req_10237_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2645), ack => type_cast_749_inst_req_0); -- 
    -- CP-element group 2646 transition  input  output  no-bypass 
    -- predecessors 2645 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_743/$exit
      -- 
    ack_10238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_749_inst_ack_0, ack => cp_elements(2646)); -- 
    phi_stmt_743_req_10239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2646), ack => phi_stmt_743_req_1); -- 
    -- CP-element group 2647 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2648 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/$entry
      -- 
    cp_elements(2647) <= cp_elements(2644);
    req_10249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2647), ack => type_cast_756_inst_req_0); -- 
    -- CP-element group 2648 transition  input  output  no-bypass 
    -- predecessors 2647 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_750/$exit
      -- 
    ack_10250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_756_inst_ack_0, ack => cp_elements(2648)); -- 
    phi_stmt_750_req_10251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2648), ack => phi_stmt_750_req_1); -- 
    -- CP-element group 2649 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2650 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/$entry
      -- 
    cp_elements(2649) <= cp_elements(2644);
    req_10261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2649), ack => type_cast_763_inst_req_0); -- 
    -- CP-element group 2650 transition  input  output  no-bypass 
    -- predecessors 2649 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_757/$exit
      -- 
    ack_10262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_0, ack => cp_elements(2650)); -- 
    phi_stmt_757_req_10263_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2650), ack => phi_stmt_757_req_1); -- 
    -- CP-element group 2651 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2652 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/$entry
      -- 
    cp_elements(2651) <= cp_elements(2644);
    req_10273_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2651), ack => type_cast_770_inst_req_0); -- 
    -- CP-element group 2652 transition  input  output  no-bypass 
    -- predecessors 2651 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_764/$exit
      -- 
    ack_10274_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_770_inst_ack_0, ack => cp_elements(2652)); -- 
    phi_stmt_764_req_10275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2652), ack => phi_stmt_764_req_1); -- 
    -- CP-element group 2653 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2654 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/$entry
      -- 
    cp_elements(2653) <= cp_elements(2644);
    req_10285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2653), ack => type_cast_777_inst_req_0); -- 
    -- CP-element group 2654 transition  input  output  no-bypass 
    -- predecessors 2653 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_771/$exit
      -- 
    ack_10286_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_777_inst_ack_0, ack => cp_elements(2654)); -- 
    phi_stmt_771_req_10287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2654), ack => phi_stmt_771_req_1); -- 
    -- CP-element group 2655 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2656 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/req
      -- 
    cp_elements(2655) <= cp_elements(2644);
    req_10297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2655), ack => type_cast_784_inst_req_0); -- 
    -- CP-element group 2656 transition  input  output  no-bypass 
    -- predecessors 2655 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_req
      -- 
    ack_10298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_0, ack => cp_elements(2656)); -- 
    phi_stmt_778_req_10299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2656), ack => phi_stmt_778_req_1); -- 
    -- CP-element group 2657 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2658 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/req
      -- 
    cp_elements(2657) <= cp_elements(2644);
    req_10309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2657), ack => type_cast_791_inst_req_0); -- 
    -- CP-element group 2658 transition  input  output  no-bypass 
    -- predecessors 2657 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_req
      -- 
    ack_10310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_791_inst_ack_0, ack => cp_elements(2658)); -- 
    phi_stmt_785_req_10311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2658), ack => phi_stmt_785_req_1); -- 
    -- CP-element group 2659 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2660 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/req
      -- 
    cp_elements(2659) <= cp_elements(2644);
    req_10321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2659), ack => type_cast_798_inst_req_0); -- 
    -- CP-element group 2660 transition  input  output  no-bypass 
    -- predecessors 2659 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_req
      -- 
    ack_10322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_798_inst_ack_0, ack => cp_elements(2660)); -- 
    phi_stmt_792_req_10323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2660), ack => phi_stmt_792_req_1); -- 
    -- CP-element group 2661 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2662 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/req
      -- 
    cp_elements(2661) <= cp_elements(2644);
    req_10333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2661), ack => type_cast_805_inst_req_0); -- 
    -- CP-element group 2662 transition  input  output  no-bypass 
    -- predecessors 2661 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/ack
      -- 
    ack_10334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_805_inst_ack_0, ack => cp_elements(2662)); -- 
    phi_stmt_799_req_10335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2662), ack => phi_stmt_799_req_1); -- 
    -- CP-element group 2663 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2664 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/$entry
      -- 
    cp_elements(2663) <= cp_elements(2644);
    req_10345_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2663), ack => type_cast_812_inst_req_0); -- 
    -- CP-element group 2664 transition  input  output  no-bypass 
    -- predecessors 2663 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_806/$exit
      -- 
    ack_10346_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_812_inst_ack_0, ack => cp_elements(2664)); -- 
    phi_stmt_806_req_10347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2664), ack => phi_stmt_806_req_1); -- 
    -- CP-element group 2665 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2666 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/$entry
      -- 
    cp_elements(2665) <= cp_elements(2644);
    req_10357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2665), ack => type_cast_819_inst_req_0); -- 
    -- CP-element group 2666 transition  input  output  no-bypass 
    -- predecessors 2665 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_813/$exit
      -- 
    ack_10358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_819_inst_ack_0, ack => cp_elements(2666)); -- 
    phi_stmt_813_req_10359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2666), ack => phi_stmt_813_req_1); -- 
    -- CP-element group 2667 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2668 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/req
      -- 
    cp_elements(2667) <= cp_elements(2644);
    req_10369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2667), ack => type_cast_826_inst_req_0); -- 
    -- CP-element group 2668 transition  input  output  no-bypass 
    -- predecessors 2667 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_req
      -- 
    ack_10370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_826_inst_ack_0, ack => cp_elements(2668)); -- 
    phi_stmt_820_req_10371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2668), ack => phi_stmt_820_req_1); -- 
    -- CP-element group 2669 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2670 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/req
      -- 
    cp_elements(2669) <= cp_elements(2644);
    req_10381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2669), ack => type_cast_833_inst_req_0); -- 
    -- CP-element group 2670 transition  input  output  no-bypass 
    -- predecessors 2669 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_req
      -- 
    ack_10382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_0, ack => cp_elements(2670)); -- 
    phi_stmt_827_req_10383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2670), ack => phi_stmt_827_req_1); -- 
    -- CP-element group 2671 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2672 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/req
      -- 
    cp_elements(2671) <= cp_elements(2644);
    req_10393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2671), ack => type_cast_840_inst_req_0); -- 
    -- CP-element group 2672 transition  input  output  no-bypass 
    -- predecessors 2671 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_req
      -- 
    ack_10394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_840_inst_ack_0, ack => cp_elements(2672)); -- 
    phi_stmt_834_req_10395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2672), ack => phi_stmt_834_req_1); -- 
    -- CP-element group 2673 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2674 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/$entry
      -- 
    cp_elements(2673) <= cp_elements(2644);
    req_10405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2673), ack => type_cast_847_inst_req_0); -- 
    -- CP-element group 2674 transition  input  output  no-bypass 
    -- predecessors 2673 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_841/$exit
      -- 
    ack_10406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_0, ack => cp_elements(2674)); -- 
    phi_stmt_841_req_10407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2674), ack => phi_stmt_841_req_1); -- 
    -- CP-element group 2675 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2676 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/$entry
      -- 
    cp_elements(2675) <= cp_elements(2644);
    req_10417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2675), ack => type_cast_854_inst_req_0); -- 
    -- CP-element group 2676 transition  input  output  no-bypass 
    -- predecessors 2675 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_req
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_848/$exit
      -- 
    ack_10418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => cp_elements(2676)); -- 
    phi_stmt_848_req_10419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2676), ack => phi_stmt_848_req_1); -- 
    -- CP-element group 2677 transition  output  bypass 
    -- predecessors 2644 
    -- successors 2678 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/$entry
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/req
      -- 
    cp_elements(2677) <= cp_elements(2644);
    req_10429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2677), ack => type_cast_861_inst_req_0); -- 
    -- CP-element group 2678 transition  input  output  no-bypass 
    -- predecessors 2677 
    -- successors 2679 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/$exit
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/ack
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_req
      -- 
    ack_10430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_0, ack => cp_elements(2678)); -- 
    phi_stmt_855_req_10431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2678), ack => phi_stmt_855_req_1); -- 
    -- CP-element group 2679 join  transition  bypass 
    -- predecessors 2646 2648 2650 2652 2654 2656 2658 2660 2662 2664 2666 2668 2670 2672 2674 2676 2678 
    -- successors 2699 
    -- members (1) 
      -- 	branch_block_stmt_552/bb_3_bb_3_PhiReq/$exit
      -- 
    cpelement_group_2679 : Block -- 
      signal predecessors: BooleanArray(16 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2646);
      predecessors(1) <= cp_elements(2648);
      predecessors(2) <= cp_elements(2650);
      predecessors(3) <= cp_elements(2652);
      predecessors(4) <= cp_elements(2654);
      predecessors(5) <= cp_elements(2656);
      predecessors(6) <= cp_elements(2658);
      predecessors(7) <= cp_elements(2660);
      predecessors(8) <= cp_elements(2662);
      predecessors(9) <= cp_elements(2664);
      predecessors(10) <= cp_elements(2666);
      predecessors(11) <= cp_elements(2668);
      predecessors(12) <= cp_elements(2670);
      predecessors(13) <= cp_elements(2672);
      predecessors(14) <= cp_elements(2674);
      predecessors(15) <= cp_elements(2676);
      predecessors(16) <= cp_elements(2678);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2679)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2679),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2680 fork  transition  bypass 
    -- predecessors 2 
    -- successors 2681 2682 2683 2684 2685 2686 2687 2688 2689 2690 2691 2692 2693 2694 2695 2696 2697 
    -- members (1) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/$entry
      -- 
    cp_elements(2680) <= cp_elements(2);
    -- CP-element group 2681 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_743/phi_stmt_743_sources/type_cast_749/req
      -- 
    cp_elements(2681) <= cp_elements(2680);
    phi_stmt_743_req_10446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2681), ack => phi_stmt_743_req_0); -- 
    -- CP-element group 2682 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_750/phi_stmt_750_sources/type_cast_756/$entry
      -- 
    cp_elements(2682) <= cp_elements(2680);
    phi_stmt_750_req_10458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2682), ack => phi_stmt_750_req_0); -- 
    -- CP-element group 2683 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_757/phi_stmt_757_sources/type_cast_763/$exit
      -- 
    cp_elements(2683) <= cp_elements(2680);
    phi_stmt_757_req_10470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2683), ack => phi_stmt_757_req_0); -- 
    -- CP-element group 2684 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/type_cast_770/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/phi_stmt_764_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_764/$entry
      -- 
    cp_elements(2684) <= cp_elements(2680);
    phi_stmt_764_req_10482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2684), ack => phi_stmt_764_req_0); -- 
    -- CP-element group 2685 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/type_cast_777/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_771/phi_stmt_771_sources/$exit
      -- 
    cp_elements(2685) <= cp_elements(2680);
    phi_stmt_771_req_10494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2685), ack => phi_stmt_771_req_0); -- 
    -- CP-element group 2686 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/phi_stmt_778_sources/type_cast_784/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_778/$entry
      -- 
    cp_elements(2686) <= cp_elements(2680);
    phi_stmt_778_req_10506_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2686), ack => phi_stmt_778_req_0); -- 
    -- CP-element group 2687 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_sources/type_cast_791/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_785/phi_stmt_785_req
      -- 
    cp_elements(2687) <= cp_elements(2680);
    phi_stmt_785_req_10518_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2687), ack => phi_stmt_785_req_0); -- 
    -- CP-element group 2688 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/phi_stmt_792_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_792/$exit
      -- 
    cp_elements(2688) <= cp_elements(2680);
    phi_stmt_792_req_10530_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2688), ack => phi_stmt_792_req_0); -- 
    -- CP-element group 2689 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_799/phi_stmt_799_sources/type_cast_805/$entry
      -- 
    cp_elements(2689) <= cp_elements(2680);
    phi_stmt_799_req_10542_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2689), ack => phi_stmt_799_req_0); -- 
    -- CP-element group 2690 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_806/phi_stmt_806_sources/type_cast_812/$exit
      -- 
    cp_elements(2690) <= cp_elements(2680);
    phi_stmt_806_req_10554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2690), ack => phi_stmt_806_req_0); -- 
    -- CP-element group 2691 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/type_cast_819/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_813/phi_stmt_813_req
      -- 
    cp_elements(2691) <= cp_elements(2680);
    phi_stmt_813_req_10566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2691), ack => phi_stmt_813_req_0); -- 
    -- CP-element group 2692 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_sources/type_cast_826/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_820/phi_stmt_820_req
      -- 
    cp_elements(2692) <= cp_elements(2680);
    phi_stmt_820_req_10578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2692), ack => phi_stmt_820_req_0); -- 
    -- CP-element group 2693 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_sources/type_cast_833/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_827/phi_stmt_827_req
      -- 
    cp_elements(2693) <= cp_elements(2680);
    phi_stmt_827_req_10590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2693), ack => phi_stmt_827_req_0); -- 
    -- CP-element group 2694 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_sources/type_cast_840/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_834/phi_stmt_834_req
      -- 
    cp_elements(2694) <= cp_elements(2680);
    phi_stmt_834_req_10602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2694), ack => phi_stmt_834_req_0); -- 
    -- CP-element group 2695 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_sources/type_cast_847/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_841/phi_stmt_841_req
      -- 
    cp_elements(2695) <= cp_elements(2680);
    phi_stmt_841_req_10614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2695), ack => phi_stmt_841_req_0); -- 
    -- CP-element group 2696 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_sources/type_cast_854/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_848/phi_stmt_848_req
      -- 
    cp_elements(2696) <= cp_elements(2680);
    phi_stmt_848_req_10626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2696), ack => phi_stmt_848_req_0); -- 
    -- CP-element group 2697 transition  output  bypass 
    -- predecessors 2680 
    -- successors 2698 
    -- members (9) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/$entry
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/$exit
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/req
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_sources/type_cast_861/ack
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/phi_stmt_855/phi_stmt_855_req
      -- 
    cp_elements(2697) <= cp_elements(2680);
    phi_stmt_855_req_10638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2697), ack => phi_stmt_855_req_0); -- 
    -- CP-element group 2698 join  transition  no-bypass 
    -- predecessors 2681 2682 2683 2684 2685 2686 2687 2688 2689 2690 2691 2692 2693 2694 2695 2696 2697 
    -- successors 2699 
    -- members (1) 
      -- 	branch_block_stmt_552/bbx_xnph_bb_3_PhiReq/$exit
      -- 
    cpelement_group_2698 : Block -- 
      signal predecessors: BooleanArray(16 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2681);
      predecessors(1) <= cp_elements(2682);
      predecessors(2) <= cp_elements(2683);
      predecessors(3) <= cp_elements(2684);
      predecessors(4) <= cp_elements(2685);
      predecessors(5) <= cp_elements(2686);
      predecessors(6) <= cp_elements(2687);
      predecessors(7) <= cp_elements(2688);
      predecessors(8) <= cp_elements(2689);
      predecessors(9) <= cp_elements(2690);
      predecessors(10) <= cp_elements(2691);
      predecessors(11) <= cp_elements(2692);
      predecessors(12) <= cp_elements(2693);
      predecessors(13) <= cp_elements(2694);
      predecessors(14) <= cp_elements(2695);
      predecessors(15) <= cp_elements(2696);
      predecessors(16) <= cp_elements(2697);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(2698)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2698),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2699 merge  place  bypass 
    -- predecessors 2679 2698 
    -- successors 2700 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiReqMerge
      -- 
    cp_elements(2699) <= OrReduce(cp_elements(2679) & cp_elements(2698));
    -- CP-element group 2700 fork  transition  bypass 
    -- predecessors 2699 
    -- successors 2701 2702 2703 2704 2705 2706 2707 2708 2709 2710 2711 2712 2713 2714 2715 2716 2717 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/$entry
      -- 
    cp_elements(2700) <= cp_elements(2699);
    -- CP-element group 2701 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_743_ack
      -- 
    phi_stmt_743_ack_10643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_743_ack_0, ack => cp_elements(2701)); -- 
    -- CP-element group 2702 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_750_ack
      -- 
    phi_stmt_750_ack_10644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_750_ack_0, ack => cp_elements(2702)); -- 
    -- CP-element group 2703 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_757_ack
      -- 
    phi_stmt_757_ack_10645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_757_ack_0, ack => cp_elements(2703)); -- 
    -- CP-element group 2704 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_764_ack
      -- 
    phi_stmt_764_ack_10646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_764_ack_0, ack => cp_elements(2704)); -- 
    -- CP-element group 2705 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_771_ack
      -- 
    phi_stmt_771_ack_10647_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_771_ack_0, ack => cp_elements(2705)); -- 
    -- CP-element group 2706 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_778_ack
      -- 
    phi_stmt_778_ack_10648_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_778_ack_0, ack => cp_elements(2706)); -- 
    -- CP-element group 2707 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_785_ack
      -- 
    phi_stmt_785_ack_10649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_785_ack_0, ack => cp_elements(2707)); -- 
    -- CP-element group 2708 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_792_ack
      -- 
    phi_stmt_792_ack_10650_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_792_ack_0, ack => cp_elements(2708)); -- 
    -- CP-element group 2709 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_799_ack
      -- 
    phi_stmt_799_ack_10651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_799_ack_0, ack => cp_elements(2709)); -- 
    -- CP-element group 2710 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_806_ack
      -- 
    phi_stmt_806_ack_10652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_806_ack_0, ack => cp_elements(2710)); -- 
    -- CP-element group 2711 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_813_ack
      -- 
    phi_stmt_813_ack_10653_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_813_ack_0, ack => cp_elements(2711)); -- 
    -- CP-element group 2712 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_820_ack
      -- 
    phi_stmt_820_ack_10654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_820_ack_0, ack => cp_elements(2712)); -- 
    -- CP-element group 2713 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_827_ack
      -- 
    phi_stmt_827_ack_10655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_827_ack_0, ack => cp_elements(2713)); -- 
    -- CP-element group 2714 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_834_ack
      -- 
    phi_stmt_834_ack_10656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_834_ack_0, ack => cp_elements(2714)); -- 
    -- CP-element group 2715 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_841_ack
      -- 
    phi_stmt_841_ack_10657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_841_ack_0, ack => cp_elements(2715)); -- 
    -- CP-element group 2716 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_848_ack
      -- 
    phi_stmt_848_ack_10658_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_848_ack_0, ack => cp_elements(2716)); -- 
    -- CP-element group 2717 transition  input  no-bypass 
    -- predecessors 2700 
    -- successors 2718 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/phi_stmt_855_ack
      -- 
    phi_stmt_855_ack_10659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_855_ack_0, ack => cp_elements(2717)); -- 
    -- CP-element group 2718 join  transition  bypass 
    -- predecessors 2701 2702 2703 2704 2705 2706 2707 2708 2709 2710 2711 2712 2713 2714 2715 2716 2717 
    -- successors 3 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_742_PhiAck/$exit
      -- 
    cpelement_group_2718 : Block -- 
      signal predecessors: BooleanArray(16 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2701);
      predecessors(1) <= cp_elements(2702);
      predecessors(2) <= cp_elements(2703);
      predecessors(3) <= cp_elements(2704);
      predecessors(4) <= cp_elements(2705);
      predecessors(5) <= cp_elements(2706);
      predecessors(6) <= cp_elements(2707);
      predecessors(7) <= cp_elements(2708);
      predecessors(8) <= cp_elements(2709);
      predecessors(9) <= cp_elements(2710);
      predecessors(10) <= cp_elements(2711);
      predecessors(11) <= cp_elements(2712);
      predecessors(12) <= cp_elements(2713);
      predecessors(13) <= cp_elements(2714);
      predecessors(14) <= cp_elements(2715);
      predecessors(15) <= cp_elements(2716);
      predecessors(16) <= cp_elements(2717);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2718)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2718),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2719 transition  dead  bypass 
    -- predecessors 2344 
    -- successors 2720 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_dead_link/dead_transition
      -- 
    cp_elements(2719) <= false;
    -- CP-element group 2720 transition  bypass 
    -- predecessors 2719 
    -- successors 5 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_dead_link/$exit
      -- 
    cp_elements(2720) <= cp_elements(2719);
    -- CP-element group 2721 fork  transition  bypass 
    -- predecessors 2348 
    -- successors 2722 2724 2726 2728 2730 2732 2734 2736 2738 2740 2742 2744 2746 2748 2750 2752 
    -- members (1) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/$entry
      -- 
    cp_elements(2721) <= cp_elements(2348);
    -- CP-element group 2722 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2723 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/phi_stmt_1890_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/phi_stmt_1890_sources/type_cast_1893/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/phi_stmt_1890_sources/type_cast_1893/req
      -- 
    cp_elements(2722) <= cp_elements(2721);
    req_10676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2722), ack => type_cast_1893_inst_req_0); -- 
    -- CP-element group 2723 transition  input  output  no-bypass 
    -- predecessors 2722 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/phi_stmt_1890_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/phi_stmt_1890_sources/type_cast_1893/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/phi_stmt_1890_sources/type_cast_1893/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1890/phi_stmt_1890_req
      -- 
    ack_10677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1893_inst_ack_0, ack => cp_elements(2723)); -- 
    phi_stmt_1890_req_10678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2723), ack => phi_stmt_1890_req_0); -- 
    -- CP-element group 2724 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2725 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/phi_stmt_1894_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/phi_stmt_1894_sources/type_cast_1897/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/phi_stmt_1894_sources/type_cast_1897/req
      -- 
    cp_elements(2724) <= cp_elements(2721);
    req_10688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2724), ack => type_cast_1897_inst_req_0); -- 
    -- CP-element group 2725 transition  input  output  no-bypass 
    -- predecessors 2724 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/phi_stmt_1894_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/phi_stmt_1894_sources/type_cast_1897/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/phi_stmt_1894_sources/type_cast_1897/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1894/phi_stmt_1894_req
      -- 
    ack_10689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1897_inst_ack_0, ack => cp_elements(2725)); -- 
    phi_stmt_1894_req_10690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2725), ack => phi_stmt_1894_req_0); -- 
    -- CP-element group 2726 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2727 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/phi_stmt_1898_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/phi_stmt_1898_sources/type_cast_1901/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/phi_stmt_1898_sources/type_cast_1901/req
      -- 
    cp_elements(2726) <= cp_elements(2721);
    req_10700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2726), ack => type_cast_1901_inst_req_0); -- 
    -- CP-element group 2727 transition  input  output  no-bypass 
    -- predecessors 2726 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/phi_stmt_1898_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/phi_stmt_1898_sources/type_cast_1901/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/phi_stmt_1898_sources/type_cast_1901/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1898/phi_stmt_1898_req
      -- 
    ack_10701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1901_inst_ack_0, ack => cp_elements(2727)); -- 
    phi_stmt_1898_req_10702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2727), ack => phi_stmt_1898_req_0); -- 
    -- CP-element group 2728 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2729 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/phi_stmt_1902_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/phi_stmt_1902_sources/type_cast_1905/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/phi_stmt_1902_sources/type_cast_1905/req
      -- 
    cp_elements(2728) <= cp_elements(2721);
    req_10712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2728), ack => type_cast_1905_inst_req_0); -- 
    -- CP-element group 2729 transition  input  output  no-bypass 
    -- predecessors 2728 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/phi_stmt_1902_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/phi_stmt_1902_sources/type_cast_1905/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/phi_stmt_1902_sources/type_cast_1905/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1902/phi_stmt_1902_req
      -- 
    ack_10713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1905_inst_ack_0, ack => cp_elements(2729)); -- 
    phi_stmt_1902_req_10714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2729), ack => phi_stmt_1902_req_0); -- 
    -- CP-element group 2730 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2731 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/phi_stmt_1906_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/phi_stmt_1906_sources/type_cast_1909/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/phi_stmt_1906_sources/type_cast_1909/req
      -- 
    cp_elements(2730) <= cp_elements(2721);
    req_10724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2730), ack => type_cast_1909_inst_req_0); -- 
    -- CP-element group 2731 transition  input  output  no-bypass 
    -- predecessors 2730 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/phi_stmt_1906_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/phi_stmt_1906_sources/type_cast_1909/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/phi_stmt_1906_sources/type_cast_1909/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1906/phi_stmt_1906_req
      -- 
    ack_10725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1909_inst_ack_0, ack => cp_elements(2731)); -- 
    phi_stmt_1906_req_10726_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2731), ack => phi_stmt_1906_req_0); -- 
    -- CP-element group 2732 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2733 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1913/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1913/req
      -- 
    cp_elements(2732) <= cp_elements(2721);
    req_10736_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2732), ack => type_cast_1913_inst_req_0); -- 
    -- CP-element group 2733 transition  input  output  no-bypass 
    -- predecessors 2732 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1913/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1913/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1910/phi_stmt_1910_req
      -- 
    ack_10737_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1913_inst_ack_0, ack => cp_elements(2733)); -- 
    phi_stmt_1910_req_10738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2733), ack => phi_stmt_1910_req_0); -- 
    -- CP-element group 2734 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2735 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/req
      -- 
    cp_elements(2734) <= cp_elements(2721);
    req_10748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2734), ack => type_cast_1917_inst_req_0); -- 
    -- CP-element group 2735 transition  input  output  no-bypass 
    -- predecessors 2734 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/phi_stmt_1914_sources/type_cast_1917/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1914/phi_stmt_1914_req
      -- 
    ack_10749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1917_inst_ack_0, ack => cp_elements(2735)); -- 
    phi_stmt_1914_req_10750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2735), ack => phi_stmt_1914_req_0); -- 
    -- CP-element group 2736 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2737 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/phi_stmt_1918_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/phi_stmt_1918_sources/type_cast_1921/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/phi_stmt_1918_sources/type_cast_1921/req
      -- 
    cp_elements(2736) <= cp_elements(2721);
    req_10760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2736), ack => type_cast_1921_inst_req_0); -- 
    -- CP-element group 2737 transition  input  output  no-bypass 
    -- predecessors 2736 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/phi_stmt_1918_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/phi_stmt_1918_sources/type_cast_1921/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/phi_stmt_1918_sources/type_cast_1921/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1918/phi_stmt_1918_req
      -- 
    ack_10761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1921_inst_ack_0, ack => cp_elements(2737)); -- 
    phi_stmt_1918_req_10762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2737), ack => phi_stmt_1918_req_0); -- 
    -- CP-element group 2738 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2739 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/phi_stmt_1922_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/phi_stmt_1922_sources/type_cast_1925/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/phi_stmt_1922_sources/type_cast_1925/req
      -- 
    cp_elements(2738) <= cp_elements(2721);
    req_10772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2738), ack => type_cast_1925_inst_req_0); -- 
    -- CP-element group 2739 transition  input  output  no-bypass 
    -- predecessors 2738 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/phi_stmt_1922_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/phi_stmt_1922_sources/type_cast_1925/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/phi_stmt_1922_sources/type_cast_1925/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1922/phi_stmt_1922_req
      -- 
    ack_10773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1925_inst_ack_0, ack => cp_elements(2739)); -- 
    phi_stmt_1922_req_10774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2739), ack => phi_stmt_1922_req_0); -- 
    -- CP-element group 2740 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2741 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/phi_stmt_1926_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/phi_stmt_1926_sources/type_cast_1929/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/phi_stmt_1926_sources/type_cast_1929/req
      -- 
    cp_elements(2740) <= cp_elements(2721);
    req_10784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2740), ack => type_cast_1929_inst_req_0); -- 
    -- CP-element group 2741 transition  input  output  no-bypass 
    -- predecessors 2740 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/phi_stmt_1926_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/phi_stmt_1926_sources/type_cast_1929/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/phi_stmt_1926_sources/type_cast_1929/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1926/phi_stmt_1926_req
      -- 
    ack_10785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1929_inst_ack_0, ack => cp_elements(2741)); -- 
    phi_stmt_1926_req_10786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2741), ack => phi_stmt_1926_req_0); -- 
    -- CP-element group 2742 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2743 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/phi_stmt_1930_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/phi_stmt_1930_sources/type_cast_1933/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/phi_stmt_1930_sources/type_cast_1933/req
      -- 
    cp_elements(2742) <= cp_elements(2721);
    req_10796_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2742), ack => type_cast_1933_inst_req_0); -- 
    -- CP-element group 2743 transition  input  output  no-bypass 
    -- predecessors 2742 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/phi_stmt_1930_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/phi_stmt_1930_sources/type_cast_1933/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/phi_stmt_1930_sources/type_cast_1933/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1930/phi_stmt_1930_req
      -- 
    ack_10797_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1933_inst_ack_0, ack => cp_elements(2743)); -- 
    phi_stmt_1930_req_10798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2743), ack => phi_stmt_1930_req_0); -- 
    -- CP-element group 2744 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2745 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/req
      -- 
    cp_elements(2744) <= cp_elements(2721);
    req_10808_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2744), ack => type_cast_1937_inst_req_0); -- 
    -- CP-element group 2745 transition  input  output  no-bypass 
    -- predecessors 2744 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/phi_stmt_1934_sources/type_cast_1937/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1934/phi_stmt_1934_req
      -- 
    ack_10809_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1937_inst_ack_0, ack => cp_elements(2745)); -- 
    phi_stmt_1934_req_10810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2745), ack => phi_stmt_1934_req_0); -- 
    -- CP-element group 2746 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2747 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/phi_stmt_1938_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/phi_stmt_1938_sources/type_cast_1941/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/phi_stmt_1938_sources/type_cast_1941/req
      -- 
    cp_elements(2746) <= cp_elements(2721);
    req_10820_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2746), ack => type_cast_1941_inst_req_0); -- 
    -- CP-element group 2747 transition  input  output  no-bypass 
    -- predecessors 2746 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/phi_stmt_1938_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/phi_stmt_1938_sources/type_cast_1941/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/phi_stmt_1938_sources/type_cast_1941/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1938/phi_stmt_1938_req
      -- 
    ack_10821_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_0, ack => cp_elements(2747)); -- 
    phi_stmt_1938_req_10822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2747), ack => phi_stmt_1938_req_0); -- 
    -- CP-element group 2748 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2749 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/phi_stmt_1942_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/phi_stmt_1942_sources/type_cast_1945/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/phi_stmt_1942_sources/type_cast_1945/req
      -- 
    cp_elements(2748) <= cp_elements(2721);
    req_10832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2748), ack => type_cast_1945_inst_req_0); -- 
    -- CP-element group 2749 transition  input  output  no-bypass 
    -- predecessors 2748 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/phi_stmt_1942_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/phi_stmt_1942_sources/type_cast_1945/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/phi_stmt_1942_sources/type_cast_1945/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1942/phi_stmt_1942_req
      -- 
    ack_10833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1945_inst_ack_0, ack => cp_elements(2749)); -- 
    phi_stmt_1942_req_10834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2749), ack => phi_stmt_1942_req_0); -- 
    -- CP-element group 2750 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2751 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/phi_stmt_1946_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/phi_stmt_1946_sources/type_cast_1949/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/phi_stmt_1946_sources/type_cast_1949/req
      -- 
    cp_elements(2750) <= cp_elements(2721);
    req_10844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2750), ack => type_cast_1949_inst_req_0); -- 
    -- CP-element group 2751 transition  input  output  no-bypass 
    -- predecessors 2750 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/phi_stmt_1946_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/phi_stmt_1946_sources/type_cast_1949/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/phi_stmt_1946_sources/type_cast_1949/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1946/phi_stmt_1946_req
      -- 
    ack_10845_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1949_inst_ack_0, ack => cp_elements(2751)); -- 
    phi_stmt_1946_req_10846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2751), ack => phi_stmt_1946_req_0); -- 
    -- CP-element group 2752 transition  output  bypass 
    -- predecessors 2721 
    -- successors 2753 
    -- members (4) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/phi_stmt_1950_sources/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/phi_stmt_1950_sources/type_cast_1953/$entry
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/phi_stmt_1950_sources/type_cast_1953/req
      -- 
    cp_elements(2752) <= cp_elements(2721);
    req_10856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2752), ack => type_cast_1953_inst_req_0); -- 
    -- CP-element group 2753 transition  input  output  no-bypass 
    -- predecessors 2752 
    -- successors 2754 
    -- members (5) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/phi_stmt_1950_sources/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/phi_stmt_1950_sources/type_cast_1953/$exit
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/phi_stmt_1950_sources/type_cast_1953/ack
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/phi_stmt_1950/phi_stmt_1950_req
      -- 
    ack_10857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1953_inst_ack_0, ack => cp_elements(2753)); -- 
    phi_stmt_1950_req_10858_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2753), ack => phi_stmt_1950_req_0); -- 
    -- CP-element group 2754 join  transition  bypass 
    -- predecessors 2723 2725 2727 2729 2731 2733 2735 2737 2739 2741 2743 2745 2747 2749 2751 2753 
    -- successors 2755 
    -- members (1) 
      -- 	branch_block_stmt_552/bb_3_xx_x_crit_edge_PhiReq/$exit
      -- 
    cpelement_group_2754 : Block -- 
      signal predecessors: BooleanArray(15 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2723);
      predecessors(1) <= cp_elements(2725);
      predecessors(2) <= cp_elements(2727);
      predecessors(3) <= cp_elements(2729);
      predecessors(4) <= cp_elements(2731);
      predecessors(5) <= cp_elements(2733);
      predecessors(6) <= cp_elements(2735);
      predecessors(7) <= cp_elements(2737);
      predecessors(8) <= cp_elements(2739);
      predecessors(9) <= cp_elements(2741);
      predecessors(10) <= cp_elements(2743);
      predecessors(11) <= cp_elements(2745);
      predecessors(12) <= cp_elements(2747);
      predecessors(13) <= cp_elements(2749);
      predecessors(14) <= cp_elements(2751);
      predecessors(15) <= cp_elements(2753);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2754)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2754),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2755 place  bypass 
    -- predecessors 2754 
    -- successors 2756 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiReqMerge
      -- 
    cp_elements(2755) <= cp_elements(2754);
    -- CP-element group 2756 fork  transition  bypass 
    -- predecessors 2755 
    -- successors 2757 2758 2759 2760 2761 2762 2763 2764 2765 2766 2767 2768 2769 2770 2771 2772 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/$entry
      -- 
    cp_elements(2756) <= cp_elements(2755);
    -- CP-element group 2757 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1890_ack
      -- 
    phi_stmt_1890_ack_10863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1890_ack_0, ack => cp_elements(2757)); -- 
    -- CP-element group 2758 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1894_ack
      -- 
    phi_stmt_1894_ack_10864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1894_ack_0, ack => cp_elements(2758)); -- 
    -- CP-element group 2759 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1898_ack
      -- 
    phi_stmt_1898_ack_10865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1898_ack_0, ack => cp_elements(2759)); -- 
    -- CP-element group 2760 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1902_ack
      -- 
    phi_stmt_1902_ack_10866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1902_ack_0, ack => cp_elements(2760)); -- 
    -- CP-element group 2761 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1906_ack
      -- 
    phi_stmt_1906_ack_10867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1906_ack_0, ack => cp_elements(2761)); -- 
    -- CP-element group 2762 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1910_ack
      -- 
    phi_stmt_1910_ack_10868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1910_ack_0, ack => cp_elements(2762)); -- 
    -- CP-element group 2763 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1914_ack
      -- 
    phi_stmt_1914_ack_10869_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1914_ack_0, ack => cp_elements(2763)); -- 
    -- CP-element group 2764 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1918_ack
      -- 
    phi_stmt_1918_ack_10870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1918_ack_0, ack => cp_elements(2764)); -- 
    -- CP-element group 2765 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1922_ack
      -- 
    phi_stmt_1922_ack_10871_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1922_ack_0, ack => cp_elements(2765)); -- 
    -- CP-element group 2766 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1926_ack
      -- 
    phi_stmt_1926_ack_10872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1926_ack_0, ack => cp_elements(2766)); -- 
    -- CP-element group 2767 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1930_ack
      -- 
    phi_stmt_1930_ack_10873_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1930_ack_0, ack => cp_elements(2767)); -- 
    -- CP-element group 2768 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1934_ack
      -- 
    phi_stmt_1934_ack_10874_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1934_ack_0, ack => cp_elements(2768)); -- 
    -- CP-element group 2769 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1938_ack
      -- 
    phi_stmt_1938_ack_10875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1938_ack_0, ack => cp_elements(2769)); -- 
    -- CP-element group 2770 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1942_ack
      -- 
    phi_stmt_1942_ack_10876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1942_ack_0, ack => cp_elements(2770)); -- 
    -- CP-element group 2771 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1946_ack
      -- 
    phi_stmt_1946_ack_10877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1946_ack_0, ack => cp_elements(2771)); -- 
    -- CP-element group 2772 transition  input  no-bypass 
    -- predecessors 2756 
    -- successors 2773 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/phi_stmt_1950_ack
      -- 
    phi_stmt_1950_ack_10878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1950_ack_0, ack => cp_elements(2772)); -- 
    -- CP-element group 2773 join  transition  bypass 
    -- predecessors 2757 2758 2759 2760 2761 2762 2763 2764 2765 2766 2767 2768 2769 2770 2771 2772 
    -- successors 5 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_1889_PhiAck/$exit
      -- 
    cpelement_group_2773 : Block -- 
      signal predecessors: BooleanArray(15 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(2757);
      predecessors(1) <= cp_elements(2758);
      predecessors(2) <= cp_elements(2759);
      predecessors(3) <= cp_elements(2760);
      predecessors(4) <= cp_elements(2761);
      predecessors(5) <= cp_elements(2762);
      predecessors(6) <= cp_elements(2763);
      predecessors(7) <= cp_elements(2764);
      predecessors(8) <= cp_elements(2765);
      predecessors(9) <= cp_elements(2766);
      predecessors(10) <= cp_elements(2767);
      predecessors(11) <= cp_elements(2768);
      predecessors(12) <= cp_elements(2769);
      predecessors(13) <= cp_elements(2770);
      predecessors(14) <= cp_elements(2771);
      predecessors(15) <= cp_elements(2772);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(2773)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2773),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 2774 transition  dead  bypass 
    -- predecessors 2608 
    -- successors 2775 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_2037_dead_link/dead_transition
      -- 
    cp_elements(2774) <= false;
    -- CP-element group 2775 transition  bypass 
    -- predecessors 2774 
    -- successors 7 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_2037_dead_link/$exit
      -- 
    cp_elements(2775) <= cp_elements(2774);
    -- CP-element group 2776 transition  dead  bypass 
    -- predecessors 2629 
    -- successors 2777 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_2056_dead_link/dead_transition
      -- 
    cp_elements(2776) <= false;
    -- CP-element group 2777 transition  bypass 
    -- predecessors 2776 
    -- successors 8 
    -- members (1) 
      -- 	branch_block_stmt_552/merge_stmt_2056_dead_link/$exit
      -- 
    cp_elements(2777) <= cp_elements(2776);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1010_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1010_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1010_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1010_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1010_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1010_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1022_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1022_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1022_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1022_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1022_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1022_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1028_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1028_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1028_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1028_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1028_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1028_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1034_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1034_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1034_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1034_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1034_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1034_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1040_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1040_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1040_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1040_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1040_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1040_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1046_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1046_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1046_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1046_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1046_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1046_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1052_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1052_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1052_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1052_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1052_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1052_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1058_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1058_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1058_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1058_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1058_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1058_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1064_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1064_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1064_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1064_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1064_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1064_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1070_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1070_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1070_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1070_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1070_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1070_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1076_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1076_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1076_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1076_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1076_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1076_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1082_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1082_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1082_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1082_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1082_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1082_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1088_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1088_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1088_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1088_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1088_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1088_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1094_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1094_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1094_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1094_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1094_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1094_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1100_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_1100_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1100_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1100_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_1100_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_1100_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_606_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_606_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_606_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_606_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_606_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_606_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_618_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_618_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_618_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_618_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_618_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_618_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_630_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_630_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_630_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_630_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_630_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_630_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_636_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_636_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_636_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_636_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_636_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_636_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_642_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_642_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_642_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_642_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_642_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_642_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_648_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_648_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_648_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_648_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_648_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_648_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_660_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_660_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_660_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_660_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_660_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_660_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_666_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_666_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_666_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_666_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_666_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_666_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_672_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_672_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_672_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_672_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_672_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_672_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_678_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_678_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_678_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_678_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_678_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_678_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_684_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_684_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_684_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_684_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_684_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_684_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_690_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_690_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_690_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_690_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_690_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_690_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_696_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_696_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_696_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_696_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_696_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_696_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_702_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_702_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_702_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_702_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_702_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_702_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_708_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_708_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_708_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_708_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_708_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_708_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_714_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_714_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_714_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_714_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_714_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_714_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_872_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_872_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_872_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_872_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_872_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_872_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_884_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_884_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_884_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_884_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_884_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_884_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_896_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_896_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_896_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_896_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_896_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_896_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_902_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_902_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_902_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_902_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_902_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_902_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_908_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_908_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_908_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_908_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_908_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_908_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_914_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_914_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_914_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_914_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_914_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_914_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_926_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_926_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_926_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_926_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_926_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_926_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_932_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_932_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_932_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_932_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_932_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_932_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_938_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_938_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_938_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_938_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_938_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_938_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_944_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_944_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_944_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_944_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_944_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_944_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_950_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_950_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_950_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_950_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_950_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_950_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_956_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_956_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_956_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_956_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_956_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_956_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_962_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_962_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_962_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_962_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_962_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_962_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_968_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_968_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_968_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_968_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_968_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_968_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_974_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_974_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_974_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_974_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_974_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_974_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_980_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_980_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_980_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_980_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_980_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_980_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_998_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_998_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_998_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_998_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_998_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_998_root_address : std_logic_vector(8 downto 0);
    signal exitcond222_1882 : std_logic_vector(0 downto 0);
    signal exitcond310_2049 : std_logic_vector(0 downto 0);
    signal exitcond_2030 : std_logic_vector(0 downto 0);
    signal iNsTr_100_1564 : std_logic_vector(31 downto 0);
    signal iNsTr_101_1569 : std_logic_vector(31 downto 0);
    signal iNsTr_102_1574 : std_logic_vector(31 downto 0);
    signal iNsTr_103_1579 : std_logic_vector(31 downto 0);
    signal iNsTr_104_1584 : std_logic_vector(31 downto 0);
    signal iNsTr_105_1589 : std_logic_vector(31 downto 0);
    signal iNsTr_106_1594 : std_logic_vector(31 downto 0);
    signal iNsTr_107_1599 : std_logic_vector(31 downto 0);
    signal iNsTr_108_1604 : std_logic_vector(31 downto 0);
    signal iNsTr_109_1609 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1134 : std_logic_vector(31 downto 0);
    signal iNsTr_110_1614 : std_logic_vector(31 downto 0);
    signal iNsTr_111_1619 : std_logic_vector(31 downto 0);
    signal iNsTr_112_1624 : std_logic_vector(31 downto 0);
    signal iNsTr_113_1629 : std_logic_vector(31 downto 0);
    signal iNsTr_114_1634 : std_logic_vector(31 downto 0);
    signal iNsTr_115_1639 : std_logic_vector(31 downto 0);
    signal iNsTr_116_1644 : std_logic_vector(31 downto 0);
    signal iNsTr_117_1649 : std_logic_vector(31 downto 0);
    signal iNsTr_118_1654 : std_logic_vector(31 downto 0);
    signal iNsTr_119_1659 : std_logic_vector(31 downto 0);
    signal iNsTr_11_1139 : std_logic_vector(31 downto 0);
    signal iNsTr_120_1664 : std_logic_vector(31 downto 0);
    signal iNsTr_121_1669 : std_logic_vector(31 downto 0);
    signal iNsTr_122_1674 : std_logic_vector(31 downto 0);
    signal iNsTr_123_1679 : std_logic_vector(31 downto 0);
    signal iNsTr_124_1684 : std_logic_vector(31 downto 0);
    signal iNsTr_125_1689 : std_logic_vector(31 downto 0);
    signal iNsTr_126_1694 : std_logic_vector(31 downto 0);
    signal iNsTr_127_1698 : std_logic_vector(31 downto 0);
    signal iNsTr_128_1702 : std_logic_vector(31 downto 0);
    signal iNsTr_129_1706 : std_logic_vector(31 downto 0);
    signal iNsTr_12_1144 : std_logic_vector(31 downto 0);
    signal iNsTr_130_1710 : std_logic_vector(31 downto 0);
    signal iNsTr_131_1715 : std_logic_vector(31 downto 0);
    signal iNsTr_132_1720 : std_logic_vector(31 downto 0);
    signal iNsTr_133_1725 : std_logic_vector(31 downto 0);
    signal iNsTr_134_1730 : std_logic_vector(31 downto 0);
    signal iNsTr_135_1735 : std_logic_vector(31 downto 0);
    signal iNsTr_136_1740 : std_logic_vector(31 downto 0);
    signal iNsTr_137_1745 : std_logic_vector(31 downto 0);
    signal iNsTr_138_1750 : std_logic_vector(31 downto 0);
    signal iNsTr_139_1755 : std_logic_vector(31 downto 0);
    signal iNsTr_13_1149 : std_logic_vector(31 downto 0);
    signal iNsTr_140_1760 : std_logic_vector(31 downto 0);
    signal iNsTr_141_1765 : std_logic_vector(31 downto 0);
    signal iNsTr_142_1770 : std_logic_vector(31 downto 0);
    signal iNsTr_143_1775 : std_logic_vector(31 downto 0);
    signal iNsTr_144_1780 : std_logic_vector(31 downto 0);
    signal iNsTr_145_1785 : std_logic_vector(31 downto 0);
    signal iNsTr_146_1790 : std_logic_vector(31 downto 0);
    signal iNsTr_147_1795 : std_logic_vector(31 downto 0);
    signal iNsTr_148_1800 : std_logic_vector(31 downto 0);
    signal iNsTr_149_1805 : std_logic_vector(31 downto 0);
    signal iNsTr_14_1154 : std_logic_vector(31 downto 0);
    signal iNsTr_150_1810 : std_logic_vector(31 downto 0);
    signal iNsTr_151_1815 : std_logic_vector(31 downto 0);
    signal iNsTr_152_1820 : std_logic_vector(31 downto 0);
    signal iNsTr_153_1825 : std_logic_vector(31 downto 0);
    signal iNsTr_154_1830 : std_logic_vector(31 downto 0);
    signal iNsTr_155_1835 : std_logic_vector(31 downto 0);
    signal iNsTr_156_1840 : std_logic_vector(31 downto 0);
    signal iNsTr_157_1845 : std_logic_vector(31 downto 0);
    signal iNsTr_158_1850 : std_logic_vector(31 downto 0);
    signal iNsTr_159_1855 : std_logic_vector(31 downto 0);
    signal iNsTr_15_1159 : std_logic_vector(31 downto 0);
    signal iNsTr_160_1860 : std_logic_vector(31 downto 0);
    signal iNsTr_161_1865 : std_logic_vector(31 downto 0);
    signal iNsTr_162_1870 : std_logic_vector(31 downto 0);
    signal iNsTr_16_1164 : std_logic_vector(31 downto 0);
    signal iNsTr_17_1169 : std_logic_vector(31 downto 0);
    signal iNsTr_18_1174 : std_logic_vector(31 downto 0);
    signal iNsTr_19_1178 : std_logic_vector(31 downto 0);
    signal iNsTr_20_1182 : std_logic_vector(31 downto 0);
    signal iNsTr_21_1186 : std_logic_vector(31 downto 0);
    signal iNsTr_22_1190 : std_logic_vector(31 downto 0);
    signal iNsTr_23_1195 : std_logic_vector(31 downto 0);
    signal iNsTr_24_1200 : std_logic_vector(31 downto 0);
    signal iNsTr_25_1205 : std_logic_vector(31 downto 0);
    signal iNsTr_26_1210 : std_logic_vector(31 downto 0);
    signal iNsTr_27_1215 : std_logic_vector(31 downto 0);
    signal iNsTr_28_1220 : std_logic_vector(31 downto 0);
    signal iNsTr_29_1225 : std_logic_vector(31 downto 0);
    signal iNsTr_30_1230 : std_logic_vector(31 downto 0);
    signal iNsTr_31_1234 : std_logic_vector(31 downto 0);
    signal iNsTr_32_1238 : std_logic_vector(31 downto 0);
    signal iNsTr_33_1242 : std_logic_vector(31 downto 0);
    signal iNsTr_34_1246 : std_logic_vector(31 downto 0);
    signal iNsTr_35_1251 : std_logic_vector(31 downto 0);
    signal iNsTr_36_1256 : std_logic_vector(31 downto 0);
    signal iNsTr_37_1261 : std_logic_vector(31 downto 0);
    signal iNsTr_38_1266 : std_logic_vector(31 downto 0);
    signal iNsTr_39_1271 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1106 : std_logic_vector(31 downto 0);
    signal iNsTr_40_1276 : std_logic_vector(31 downto 0);
    signal iNsTr_41_1281 : std_logic_vector(31 downto 0);
    signal iNsTr_42_1286 : std_logic_vector(31 downto 0);
    signal iNsTr_43_1290 : std_logic_vector(31 downto 0);
    signal iNsTr_44_1294 : std_logic_vector(31 downto 0);
    signal iNsTr_45_1298 : std_logic_vector(31 downto 0);
    signal iNsTr_46_1302 : std_logic_vector(31 downto 0);
    signal iNsTr_47_1307 : std_logic_vector(31 downto 0);
    signal iNsTr_48_1312 : std_logic_vector(31 downto 0);
    signal iNsTr_49_1317 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1110 : std_logic_vector(31 downto 0);
    signal iNsTr_50_1322 : std_logic_vector(31 downto 0);
    signal iNsTr_51_1327 : std_logic_vector(31 downto 0);
    signal iNsTr_52_1332 : std_logic_vector(31 downto 0);
    signal iNsTr_53_1337 : std_logic_vector(31 downto 0);
    signal iNsTr_54_1342 : std_logic_vector(31 downto 0);
    signal iNsTr_55_1346 : std_logic_vector(31 downto 0);
    signal iNsTr_56_1350 : std_logic_vector(31 downto 0);
    signal iNsTr_57_1354 : std_logic_vector(31 downto 0);
    signal iNsTr_58_1358 : std_logic_vector(31 downto 0);
    signal iNsTr_59_1363 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1114 : std_logic_vector(31 downto 0);
    signal iNsTr_60_1368 : std_logic_vector(31 downto 0);
    signal iNsTr_61_1373 : std_logic_vector(31 downto 0);
    signal iNsTr_62_1378 : std_logic_vector(31 downto 0);
    signal iNsTr_63_1383 : std_logic_vector(31 downto 0);
    signal iNsTr_64_1388 : std_logic_vector(31 downto 0);
    signal iNsTr_65_1393 : std_logic_vector(31 downto 0);
    signal iNsTr_66_1398 : std_logic_vector(31 downto 0);
    signal iNsTr_67_1403 : std_logic_vector(31 downto 0);
    signal iNsTr_68_1408 : std_logic_vector(31 downto 0);
    signal iNsTr_69_1413 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1118 : std_logic_vector(31 downto 0);
    signal iNsTr_70_1418 : std_logic_vector(31 downto 0);
    signal iNsTr_71_1423 : std_logic_vector(31 downto 0);
    signal iNsTr_72_1428 : std_logic_vector(31 downto 0);
    signal iNsTr_73_1433 : std_logic_vector(31 downto 0);
    signal iNsTr_74_1438 : std_logic_vector(31 downto 0);
    signal iNsTr_75_1443 : std_logic_vector(31 downto 0);
    signal iNsTr_76_1448 : std_logic_vector(31 downto 0);
    signal iNsTr_77_1453 : std_logic_vector(31 downto 0);
    signal iNsTr_78_1458 : std_logic_vector(31 downto 0);
    signal iNsTr_79_1463 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1122 : std_logic_vector(31 downto 0);
    signal iNsTr_80_1468 : std_logic_vector(31 downto 0);
    signal iNsTr_81_1473 : std_logic_vector(31 downto 0);
    signal iNsTr_82_1478 : std_logic_vector(31 downto 0);
    signal iNsTr_83_1483 : std_logic_vector(31 downto 0);
    signal iNsTr_84_1488 : std_logic_vector(31 downto 0);
    signal iNsTr_85_1493 : std_logic_vector(31 downto 0);
    signal iNsTr_86_1498 : std_logic_vector(31 downto 0);
    signal iNsTr_87_1503 : std_logic_vector(31 downto 0);
    signal iNsTr_88_1508 : std_logic_vector(31 downto 0);
    signal iNsTr_89_1513 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1126 : std_logic_vector(31 downto 0);
    signal iNsTr_90_1518 : std_logic_vector(31 downto 0);
    signal iNsTr_91_1522 : std_logic_vector(31 downto 0);
    signal iNsTr_92_1526 : std_logic_vector(31 downto 0);
    signal iNsTr_93_1530 : std_logic_vector(31 downto 0);
    signal iNsTr_94_1534 : std_logic_vector(31 downto 0);
    signal iNsTr_95_1539 : std_logic_vector(31 downto 0);
    signal iNsTr_96_1544 : std_logic_vector(31 downto 0);
    signal iNsTr_97_1549 : std_logic_vector(31 downto 0);
    signal iNsTr_98_1554 : std_logic_vector(31 downto 0);
    signal iNsTr_99_1559 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1130 : std_logic_vector(31 downto 0);
    signal indvar56_589 : std_logic_vector(31 downto 0);
    signal indvar60_555 : std_logic_vector(31 downto 0);
    signal indvar_743 : std_logic_vector(31 downto 0);
    signal indvarx_xnext57_2024 : std_logic_vector(31 downto 0);
    signal indvarx_xnext61_2043 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1876 : std_logic_vector(31 downto 0);
    signal ptr_deref_1105_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1105_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1105_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1105_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1105_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1109_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1109_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1109_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1109_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1109_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1113_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1113_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1113_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1113_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1113_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1117_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1117_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1117_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1117_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1117_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1121_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1121_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1121_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1121_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1121_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1125_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1125_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1125_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1125_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1125_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1129_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1129_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1129_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1129_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1129_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1133_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1133_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1133_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1133_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1133_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1177_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1177_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1177_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1177_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1177_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1181_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1181_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1181_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1181_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1181_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1185_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1185_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1185_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1185_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1185_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1189_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1189_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1189_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1189_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1189_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1233_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1233_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1233_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1233_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1233_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1237_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1237_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1237_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1237_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1237_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1241_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1241_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1241_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1241_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1241_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1245_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1245_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1245_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1245_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1245_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1289_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1289_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1289_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1289_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1289_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1293_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1293_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1293_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1293_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1293_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1297_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1297_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1297_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1297_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1297_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1301_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1301_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1301_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1301_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1301_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1345_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1345_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1345_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1345_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1345_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1349_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1349_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1349_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1349_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1349_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1353_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1353_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1353_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1353_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1353_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1357_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1357_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1357_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1357_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1357_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1521_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1521_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1521_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1521_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1521_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1525_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1525_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1525_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1525_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1525_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1529_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1529_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1529_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1529_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1529_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1533_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1533_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1697_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1697_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1697_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1697_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1697_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1701_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1701_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1701_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1701_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1701_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1705_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1705_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1705_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1705_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1705_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1709_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1709_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1709_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1709_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1709_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1956_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1956_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1956_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1956_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1956_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1956_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1960_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1960_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1960_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1960_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1960_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1960_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1964_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1964_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1964_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1964_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1964_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1964_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1968_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1968_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1968_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1968_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1968_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1968_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1972_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1972_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1972_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1972_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1972_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1972_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1976_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1976_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1976_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1976_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1976_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1976_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1980_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1980_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1980_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1980_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1980_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1980_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1984_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1984_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1984_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1984_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1984_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1984_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1988_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1988_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1988_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1988_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1988_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1988_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1992_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1992_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1992_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1992_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1992_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1992_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1996_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1996_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1996_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_1996_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1996_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_1996_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2000_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2000_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2000_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2000_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2000_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2000_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2004_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2004_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2004_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2004_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2004_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2004_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2008_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2008_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2008_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2008_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2008_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2008_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2012_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2012_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2012_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2012_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2012_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2012_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2016_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2016_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2016_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2016_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2016_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2016_word_offset_0 : std_logic_vector(8 downto 0);
    signal scevgep100_964 : std_logic_vector(31 downto 0);
    signal scevgep101_886 : std_logic_vector(31 downto 0);
    signal scevgep129_638 : std_logic_vector(31 downto 0);
    signal scevgep131_668 : std_logic_vector(31 downto 0);
    signal scevgep133_692 : std_logic_vector(31 downto 0);
    signal scevgep134_608 : std_logic_vector(31 downto 0);
    signal scevgep135_662 : std_logic_vector(31 downto 0);
    signal scevgep136_686 : std_logic_vector(31 downto 0);
    signal scevgep137_710 : std_logic_vector(31 downto 0);
    signal scevgep138_716 : std_logic_vector(31 downto 0);
    signal scevgep139_650 : std_logic_vector(31 downto 0);
    signal scevgep140_680 : std_logic_vector(31 downto 0);
    signal scevgep141_704 : std_logic_vector(31 downto 0);
    signal scevgep142_632 : std_logic_vector(31 downto 0);
    signal scevgep143_644 : std_logic_vector(31 downto 0);
    signal scevgep144_674 : std_logic_vector(31 downto 0);
    signal scevgep145_698 : std_logic_vector(31 downto 0);
    signal scevgep146_620 : std_logic_vector(31 downto 0);
    signal scevgep64_904 : std_logic_vector(31 downto 0);
    signal scevgep66_1078 : std_logic_vector(31 downto 0);
    signal scevgep68_1054 : std_logic_vector(31 downto 0);
    signal scevgep69_1030 : std_logic_vector(31 downto 0);
    signal scevgep71_934 : std_logic_vector(31 downto 0);
    signal scevgep73_958 : std_logic_vector(31 downto 0);
    signal scevgep74_874 : std_logic_vector(31 downto 0);
    signal scevgep76_1096 : std_logic_vector(31 downto 0);
    signal scevgep77_928 : std_logic_vector(31 downto 0);
    signal scevgep78_1072 : std_logic_vector(31 downto 0);
    signal scevgep79_1048 : std_logic_vector(31 downto 0);
    signal scevgep80_1024 : std_logic_vector(31 downto 0);
    signal scevgep81_952 : std_logic_vector(31 downto 0);
    signal scevgep82_976 : std_logic_vector(31 downto 0);
    signal scevgep83_982 : std_logic_vector(31 downto 0);
    signal scevgep85_1090 : std_logic_vector(31 downto 0);
    signal scevgep86_916 : std_logic_vector(31 downto 0);
    signal scevgep87_1066 : std_logic_vector(31 downto 0);
    signal scevgep88_1042 : std_logic_vector(31 downto 0);
    signal scevgep89_1012 : std_logic_vector(31 downto 0);
    signal scevgep90_946 : std_logic_vector(31 downto 0);
    signal scevgep91_970 : std_logic_vector(31 downto 0);
    signal scevgep92_898 : std_logic_vector(31 downto 0);
    signal scevgep94_1084 : std_logic_vector(31 downto 0);
    signal scevgep95_910 : std_logic_vector(31 downto 0);
    signal scevgep96_1060 : std_logic_vector(31 downto 0);
    signal scevgep97_1036 : std_logic_vector(31 downto 0);
    signal scevgep98_1000 : std_logic_vector(31 downto 0);
    signal scevgep99_940 : std_logic_vector(31 downto 0);
    signal scevgep_1102 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1008_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1008_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1009_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1009_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1020_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1020_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1021_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1021_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1026_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1026_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1027_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1027_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1032_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1032_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1033_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1033_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1038_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1038_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1039_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1039_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1044_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1044_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1045_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1045_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1050_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1050_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1051_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1051_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1056_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1056_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1057_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1057_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1062_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1062_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1063_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1063_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1068_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1068_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1069_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1069_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1074_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1074_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1075_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1075_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1080_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1080_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1081_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1081_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1086_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1086_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1087_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1087_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1092_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1092_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1093_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1093_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1098_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1098_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1099_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_1099_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_604_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_604_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_605_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_605_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_616_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_616_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_617_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_617_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_628_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_628_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_629_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_629_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_634_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_634_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_635_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_635_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_640_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_640_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_641_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_641_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_646_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_646_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_647_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_647_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_658_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_658_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_659_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_659_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_664_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_664_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_665_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_665_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_670_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_670_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_671_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_671_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_676_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_676_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_677_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_677_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_682_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_682_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_683_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_683_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_688_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_688_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_689_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_689_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_694_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_694_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_695_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_695_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_700_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_700_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_701_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_701_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_706_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_706_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_707_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_707_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_712_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_712_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_713_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_713_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_870_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_870_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_871_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_871_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_882_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_882_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_883_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_883_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_894_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_894_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_895_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_895_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_900_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_900_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_901_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_901_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_906_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_906_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_907_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_907_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_912_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_912_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_913_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_913_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_924_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_924_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_925_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_925_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_930_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_930_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_931_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_931_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_936_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_936_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_937_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_937_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_942_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_942_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_943_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_943_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_948_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_948_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_949_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_949_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_954_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_954_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_955_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_955_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_960_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_960_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_961_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_961_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_966_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_966_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_967_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_967_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_972_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_972_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_973_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_973_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_978_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_978_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_979_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_979_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_996_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_996_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_997_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_997_scaled : std_logic_vector(8 downto 0);
    signal tmp266_988 : std_logic_vector(31 downto 0);
    signal tmp267_994 : std_logic_vector(31 downto 0);
    signal tmp268_722 : std_logic_vector(31 downto 0);
    signal tmp270_1006 : std_logic_vector(31 downto 0);
    signal tmp272_1018 : std_logic_vector(31 downto 0);
    signal tmp275_728 : std_logic_vector(31 downto 0);
    signal tmp280_734 : std_logic_vector(31 downto 0);
    signal tmp285_740 : std_logic_vector(31 downto 0);
    signal tmp311_568 : std_logic_vector(31 downto 0);
    signal tmp312_602 : std_logic_vector(31 downto 0);
    signal tmp314_614 : std_logic_vector(31 downto 0);
    signal tmp316_626 : std_logic_vector(31 downto 0);
    signal tmp318_574 : std_logic_vector(31 downto 0);
    signal tmp322_656 : std_logic_vector(31 downto 0);
    signal tmp324_580 : std_logic_vector(31 downto 0);
    signal tmp329_586 : std_logic_vector(31 downto 0);
    signal tmp335_868 : std_logic_vector(31 downto 0);
    signal tmp337_880 : std_logic_vector(31 downto 0);
    signal tmp339_892 : std_logic_vector(31 downto 0);
    signal tmp344_922 : std_logic_vector(31 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1016_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1874_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1880_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1893_wire : std_logic_vector(31 downto 0);
    signal type_cast_1897_wire : std_logic_vector(31 downto 0);
    signal type_cast_1901_wire : std_logic_vector(31 downto 0);
    signal type_cast_1905_wire : std_logic_vector(31 downto 0);
    signal type_cast_1909_wire : std_logic_vector(31 downto 0);
    signal type_cast_1913_wire : std_logic_vector(31 downto 0);
    signal type_cast_1917_wire : std_logic_vector(31 downto 0);
    signal type_cast_1921_wire : std_logic_vector(31 downto 0);
    signal type_cast_1925_wire : std_logic_vector(31 downto 0);
    signal type_cast_1929_wire : std_logic_vector(31 downto 0);
    signal type_cast_1933_wire : std_logic_vector(31 downto 0);
    signal type_cast_1937_wire : std_logic_vector(31 downto 0);
    signal type_cast_1941_wire : std_logic_vector(31 downto 0);
    signal type_cast_1945_wire : std_logic_vector(31 downto 0);
    signal type_cast_1949_wire : std_logic_vector(31 downto 0);
    signal type_cast_1953_wire : std_logic_vector(31 downto 0);
    signal type_cast_2022_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2028_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2041_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2047_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_559_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_561_wire : std_logic_vector(31 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_572_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_578_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_584_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_593_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_595_wire : std_logic_vector(31 downto 0);
    signal type_cast_600_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_612_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_720_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_726_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_732_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_747_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_749_wire : std_logic_vector(31 downto 0);
    signal type_cast_754_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_756_wire : std_logic_vector(31 downto 0);
    signal type_cast_761_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_763_wire : std_logic_vector(31 downto 0);
    signal type_cast_768_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_770_wire : std_logic_vector(31 downto 0);
    signal type_cast_775_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_777_wire : std_logic_vector(31 downto 0);
    signal type_cast_782_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_784_wire : std_logic_vector(31 downto 0);
    signal type_cast_789_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_791_wire : std_logic_vector(31 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_798_wire : std_logic_vector(31 downto 0);
    signal type_cast_803_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_805_wire : std_logic_vector(31 downto 0);
    signal type_cast_810_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_812_wire : std_logic_vector(31 downto 0);
    signal type_cast_817_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_819_wire : std_logic_vector(31 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_826_wire : std_logic_vector(31 downto 0);
    signal type_cast_831_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_833_wire : std_logic_vector(31 downto 0);
    signal type_cast_838_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_840_wire : std_logic_vector(31 downto 0);
    signal type_cast_845_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_847_wire : std_logic_vector(31 downto 0);
    signal type_cast_852_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_854_wire : std_logic_vector(31 downto 0);
    signal type_cast_859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_861_wire : std_logic_vector(31 downto 0);
    signal type_cast_866_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_986_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_992_wire_constant : std_logic_vector(31 downto 0);
    signal v00x_x09_813 : std_logic_vector(31 downto 0);
    signal v01x_x08_820 : std_logic_vector(31 downto 0);
    signal v02x_x07_827 : std_logic_vector(31 downto 0);
    signal v03x_x06_834 : std_logic_vector(31 downto 0);
    signal v10x_x05_841 : std_logic_vector(31 downto 0);
    signal v11x_x04_848 : std_logic_vector(31 downto 0);
    signal v12x_x03_855 : std_logic_vector(31 downto 0);
    signal v13x_x010_806 : std_logic_vector(31 downto 0);
    signal v20x_x011_799 : std_logic_vector(31 downto 0);
    signal v21x_x012_792 : std_logic_vector(31 downto 0);
    signal v22x_x013_785 : std_logic_vector(31 downto 0);
    signal v23x_x014_778 : std_logic_vector(31 downto 0);
    signal v30x_x015_771 : std_logic_vector(31 downto 0);
    signal v31x_x016_764 : std_logic_vector(31 downto 0);
    signal v32x_x017_757 : std_logic_vector(31 downto 0);
    signal v33x_x018_750 : std_logic_vector(31 downto 0);
    signal xx_xlcssa207_1946 : std_logic_vector(31 downto 0);
    signal xx_xlcssa208_1942 : std_logic_vector(31 downto 0);
    signal xx_xlcssa209_1938 : std_logic_vector(31 downto 0);
    signal xx_xlcssa210_1934 : std_logic_vector(31 downto 0);
    signal xx_xlcssa211_1930 : std_logic_vector(31 downto 0);
    signal xx_xlcssa212_1926 : std_logic_vector(31 downto 0);
    signal xx_xlcssa213_1922 : std_logic_vector(31 downto 0);
    signal xx_xlcssa214_1918 : std_logic_vector(31 downto 0);
    signal xx_xlcssa215_1914 : std_logic_vector(31 downto 0);
    signal xx_xlcssa216_1910 : std_logic_vector(31 downto 0);
    signal xx_xlcssa217_1906 : std_logic_vector(31 downto 0);
    signal xx_xlcssa218_1902 : std_logic_vector(31 downto 0);
    signal xx_xlcssa219_1898 : std_logic_vector(31 downto 0);
    signal xx_xlcssa220_1894 : std_logic_vector(31 downto 0);
    signal xx_xlcssa221_1890 : std_logic_vector(31 downto 0);
    signal xx_xlcssa_1950 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1010_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1010_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1010_resized_base_address <= "000000000";
    array_obj_ref_1022_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1022_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1022_resized_base_address <= "000000000";
    array_obj_ref_1028_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1028_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1028_resized_base_address <= "000000000";
    array_obj_ref_1034_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1034_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1034_resized_base_address <= "000000000";
    array_obj_ref_1040_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1040_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1040_resized_base_address <= "000000000";
    array_obj_ref_1046_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1046_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1046_resized_base_address <= "000000000";
    array_obj_ref_1052_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1052_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1052_resized_base_address <= "000000000";
    array_obj_ref_1058_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1058_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1058_resized_base_address <= "000000000";
    array_obj_ref_1064_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1064_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1064_resized_base_address <= "000000000";
    array_obj_ref_1070_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1070_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1070_resized_base_address <= "000000000";
    array_obj_ref_1076_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1076_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1076_resized_base_address <= "000000000";
    array_obj_ref_1082_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1082_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1082_resized_base_address <= "000000000";
    array_obj_ref_1088_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1088_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1088_resized_base_address <= "000000000";
    array_obj_ref_1094_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1094_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1094_resized_base_address <= "000000000";
    array_obj_ref_1100_offset_scale_factor_0 <= "000010000";
    array_obj_ref_1100_offset_scale_factor_1 <= "000000001";
    array_obj_ref_1100_resized_base_address <= "000000000";
    array_obj_ref_606_offset_scale_factor_0 <= "000010000";
    array_obj_ref_606_offset_scale_factor_1 <= "000000001";
    array_obj_ref_606_resized_base_address <= "000000000";
    array_obj_ref_618_offset_scale_factor_0 <= "000010000";
    array_obj_ref_618_offset_scale_factor_1 <= "000000001";
    array_obj_ref_618_resized_base_address <= "000000000";
    array_obj_ref_630_offset_scale_factor_0 <= "000010000";
    array_obj_ref_630_offset_scale_factor_1 <= "000000001";
    array_obj_ref_630_resized_base_address <= "000000000";
    array_obj_ref_636_offset_scale_factor_0 <= "000010000";
    array_obj_ref_636_offset_scale_factor_1 <= "000000001";
    array_obj_ref_636_resized_base_address <= "000000000";
    array_obj_ref_642_offset_scale_factor_0 <= "000010000";
    array_obj_ref_642_offset_scale_factor_1 <= "000000001";
    array_obj_ref_642_resized_base_address <= "000000000";
    array_obj_ref_648_offset_scale_factor_0 <= "000010000";
    array_obj_ref_648_offset_scale_factor_1 <= "000000001";
    array_obj_ref_648_resized_base_address <= "000000000";
    array_obj_ref_660_offset_scale_factor_0 <= "000010000";
    array_obj_ref_660_offset_scale_factor_1 <= "000000001";
    array_obj_ref_660_resized_base_address <= "000000000";
    array_obj_ref_666_offset_scale_factor_0 <= "000010000";
    array_obj_ref_666_offset_scale_factor_1 <= "000000001";
    array_obj_ref_666_resized_base_address <= "000000000";
    array_obj_ref_672_offset_scale_factor_0 <= "000010000";
    array_obj_ref_672_offset_scale_factor_1 <= "000000001";
    array_obj_ref_672_resized_base_address <= "000000000";
    array_obj_ref_678_offset_scale_factor_0 <= "000010000";
    array_obj_ref_678_offset_scale_factor_1 <= "000000001";
    array_obj_ref_678_resized_base_address <= "000000000";
    array_obj_ref_684_offset_scale_factor_0 <= "000010000";
    array_obj_ref_684_offset_scale_factor_1 <= "000000001";
    array_obj_ref_684_resized_base_address <= "000000000";
    array_obj_ref_690_offset_scale_factor_0 <= "000010000";
    array_obj_ref_690_offset_scale_factor_1 <= "000000001";
    array_obj_ref_690_resized_base_address <= "000000000";
    array_obj_ref_696_offset_scale_factor_0 <= "000010000";
    array_obj_ref_696_offset_scale_factor_1 <= "000000001";
    array_obj_ref_696_resized_base_address <= "000000000";
    array_obj_ref_702_offset_scale_factor_0 <= "000010000";
    array_obj_ref_702_offset_scale_factor_1 <= "000000001";
    array_obj_ref_702_resized_base_address <= "000000000";
    array_obj_ref_708_offset_scale_factor_0 <= "000010000";
    array_obj_ref_708_offset_scale_factor_1 <= "000000001";
    array_obj_ref_708_resized_base_address <= "000000000";
    array_obj_ref_714_offset_scale_factor_0 <= "000010000";
    array_obj_ref_714_offset_scale_factor_1 <= "000000001";
    array_obj_ref_714_resized_base_address <= "000000000";
    array_obj_ref_872_offset_scale_factor_0 <= "000010000";
    array_obj_ref_872_offset_scale_factor_1 <= "000000001";
    array_obj_ref_872_resized_base_address <= "000000000";
    array_obj_ref_884_offset_scale_factor_0 <= "000010000";
    array_obj_ref_884_offset_scale_factor_1 <= "000000001";
    array_obj_ref_884_resized_base_address <= "000000000";
    array_obj_ref_896_offset_scale_factor_0 <= "000010000";
    array_obj_ref_896_offset_scale_factor_1 <= "000000001";
    array_obj_ref_896_resized_base_address <= "000000000";
    array_obj_ref_902_offset_scale_factor_0 <= "000010000";
    array_obj_ref_902_offset_scale_factor_1 <= "000000001";
    array_obj_ref_902_resized_base_address <= "000000000";
    array_obj_ref_908_offset_scale_factor_0 <= "000010000";
    array_obj_ref_908_offset_scale_factor_1 <= "000000001";
    array_obj_ref_908_resized_base_address <= "000000000";
    array_obj_ref_914_offset_scale_factor_0 <= "000010000";
    array_obj_ref_914_offset_scale_factor_1 <= "000000001";
    array_obj_ref_914_resized_base_address <= "000000000";
    array_obj_ref_926_offset_scale_factor_0 <= "000010000";
    array_obj_ref_926_offset_scale_factor_1 <= "000000001";
    array_obj_ref_926_resized_base_address <= "000000000";
    array_obj_ref_932_offset_scale_factor_0 <= "000010000";
    array_obj_ref_932_offset_scale_factor_1 <= "000000001";
    array_obj_ref_932_resized_base_address <= "000000000";
    array_obj_ref_938_offset_scale_factor_0 <= "000010000";
    array_obj_ref_938_offset_scale_factor_1 <= "000000001";
    array_obj_ref_938_resized_base_address <= "000000000";
    array_obj_ref_944_offset_scale_factor_0 <= "000010000";
    array_obj_ref_944_offset_scale_factor_1 <= "000000001";
    array_obj_ref_944_resized_base_address <= "000000000";
    array_obj_ref_950_offset_scale_factor_0 <= "000010000";
    array_obj_ref_950_offset_scale_factor_1 <= "000000001";
    array_obj_ref_950_resized_base_address <= "000000000";
    array_obj_ref_956_offset_scale_factor_0 <= "000010000";
    array_obj_ref_956_offset_scale_factor_1 <= "000000001";
    array_obj_ref_956_resized_base_address <= "000000000";
    array_obj_ref_962_offset_scale_factor_0 <= "000010000";
    array_obj_ref_962_offset_scale_factor_1 <= "000000001";
    array_obj_ref_962_resized_base_address <= "000000000";
    array_obj_ref_968_offset_scale_factor_0 <= "000010000";
    array_obj_ref_968_offset_scale_factor_1 <= "000000001";
    array_obj_ref_968_resized_base_address <= "000000000";
    array_obj_ref_974_offset_scale_factor_0 <= "000010000";
    array_obj_ref_974_offset_scale_factor_1 <= "000000001";
    array_obj_ref_974_resized_base_address <= "000000000";
    array_obj_ref_980_offset_scale_factor_0 <= "000010000";
    array_obj_ref_980_offset_scale_factor_1 <= "000000001";
    array_obj_ref_980_resized_base_address <= "000000000";
    array_obj_ref_998_offset_scale_factor_0 <= "000010000";
    array_obj_ref_998_offset_scale_factor_1 <= "000000001";
    array_obj_ref_998_resized_base_address <= "000000000";
    ptr_deref_1105_word_offset_0 <= "000000000";
    ptr_deref_1109_word_offset_0 <= "000000000";
    ptr_deref_1113_word_offset_0 <= "000000000";
    ptr_deref_1117_word_offset_0 <= "000000000";
    ptr_deref_1121_word_offset_0 <= "000000000";
    ptr_deref_1125_word_offset_0 <= "000000000";
    ptr_deref_1129_word_offset_0 <= "000000000";
    ptr_deref_1133_word_offset_0 <= "000000000";
    ptr_deref_1177_word_offset_0 <= "000000000";
    ptr_deref_1181_word_offset_0 <= "000000000";
    ptr_deref_1185_word_offset_0 <= "000000000";
    ptr_deref_1189_word_offset_0 <= "000000000";
    ptr_deref_1233_word_offset_0 <= "000000000";
    ptr_deref_1237_word_offset_0 <= "000000000";
    ptr_deref_1241_word_offset_0 <= "000000000";
    ptr_deref_1245_word_offset_0 <= "000000000";
    ptr_deref_1289_word_offset_0 <= "000000000";
    ptr_deref_1293_word_offset_0 <= "000000000";
    ptr_deref_1297_word_offset_0 <= "000000000";
    ptr_deref_1301_word_offset_0 <= "000000000";
    ptr_deref_1345_word_offset_0 <= "000000000";
    ptr_deref_1349_word_offset_0 <= "000000000";
    ptr_deref_1353_word_offset_0 <= "000000000";
    ptr_deref_1357_word_offset_0 <= "000000000";
    ptr_deref_1521_word_offset_0 <= "000000000";
    ptr_deref_1525_word_offset_0 <= "000000000";
    ptr_deref_1529_word_offset_0 <= "000000000";
    ptr_deref_1533_word_offset_0 <= "000000000";
    ptr_deref_1697_word_offset_0 <= "000000000";
    ptr_deref_1701_word_offset_0 <= "000000000";
    ptr_deref_1705_word_offset_0 <= "000000000";
    ptr_deref_1709_word_offset_0 <= "000000000";
    ptr_deref_1956_word_offset_0 <= "000000000";
    ptr_deref_1960_word_offset_0 <= "000000000";
    ptr_deref_1964_word_offset_0 <= "000000000";
    ptr_deref_1968_word_offset_0 <= "000000000";
    ptr_deref_1972_word_offset_0 <= "000000000";
    ptr_deref_1976_word_offset_0 <= "000000000";
    ptr_deref_1980_word_offset_0 <= "000000000";
    ptr_deref_1984_word_offset_0 <= "000000000";
    ptr_deref_1988_word_offset_0 <= "000000000";
    ptr_deref_1992_word_offset_0 <= "000000000";
    ptr_deref_1996_word_offset_0 <= "000000000";
    ptr_deref_2000_word_offset_0 <= "000000000";
    ptr_deref_2004_word_offset_0 <= "000000000";
    ptr_deref_2008_word_offset_0 <= "000000000";
    ptr_deref_2012_word_offset_0 <= "000000000";
    ptr_deref_2016_word_offset_0 <= "000000000";
    type_cast_1004_wire_constant <= "00000000000000000000000000000010";
    type_cast_1016_wire_constant <= "00000000000000000000000000000001";
    type_cast_1874_wire_constant <= "00000000000000000000000000000001";
    type_cast_1880_wire_constant <= "00000000000000000000000000000100";
    type_cast_2022_wire_constant <= "00000000000000000000000000000001";
    type_cast_2028_wire_constant <= "00000000000000000000000000000100";
    type_cast_2041_wire_constant <= "00000000000000000000000000000001";
    type_cast_2047_wire_constant <= "00000000000000000000000000000100";
    type_cast_559_wire_constant <= "00000000000000000000000000000000";
    type_cast_566_wire_constant <= "00000000000000000000000000000100";
    type_cast_572_wire_constant <= "00000000000000000000000000000011";
    type_cast_578_wire_constant <= "00000000000000000000000000000010";
    type_cast_584_wire_constant <= "00000000000000000000000000000001";
    type_cast_593_wire_constant <= "00000000000000000000000000000000";
    type_cast_600_wire_constant <= "00000000000000000000000000000100";
    type_cast_612_wire_constant <= "00000000000000000000000000000011";
    type_cast_624_wire_constant <= "00000000000000000000000000000010";
    type_cast_654_wire_constant <= "00000000000000000000000000000001";
    type_cast_720_wire_constant <= "00000000000000000000000000000100";
    type_cast_726_wire_constant <= "00000000000000000000000000000001";
    type_cast_732_wire_constant <= "00000000000000000000000000000010";
    type_cast_738_wire_constant <= "00000000000000000000000000000011";
    type_cast_747_wire_constant <= "00000000000000000000000000000000";
    type_cast_754_wire_constant <= "00000000000000000000000000000000";
    type_cast_761_wire_constant <= "00000000000000000000000000000000";
    type_cast_768_wire_constant <= "00000000000000000000000000000000";
    type_cast_775_wire_constant <= "00000000000000000000000000000000";
    type_cast_782_wire_constant <= "00000000000000000000000000000000";
    type_cast_789_wire_constant <= "00000000000000000000000000000000";
    type_cast_796_wire_constant <= "00000000000000000000000000000000";
    type_cast_803_wire_constant <= "00000000000000000000000000000000";
    type_cast_810_wire_constant <= "00000000000000000000000000000000";
    type_cast_817_wire_constant <= "00000000000000000000000000000000";
    type_cast_824_wire_constant <= "00000000000000000000000000000000";
    type_cast_831_wire_constant <= "00000000000000000000000000000000";
    type_cast_838_wire_constant <= "00000000000000000000000000000000";
    type_cast_845_wire_constant <= "00000000000000000000000000000000";
    type_cast_852_wire_constant <= "00000000000000000000000000000000";
    type_cast_859_wire_constant <= "00000000000000000000000000000000";
    type_cast_866_wire_constant <= "00000000000000000000000000000100";
    type_cast_878_wire_constant <= "00000000000000000000000000000011";
    type_cast_890_wire_constant <= "00000000000000000000000000000010";
    type_cast_920_wire_constant <= "00000000000000000000000000000001";
    type_cast_986_wire_constant <= "00000000000000000000000000000100";
    type_cast_992_wire_constant <= "00000000000000000000000000000011";
    phi_stmt_1890: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1893_wire;
      req(0) <= phi_stmt_1890_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1890_ack_0,
          idata => idata,
          odata => xx_xlcssa221_1890,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1890
    phi_stmt_1894: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1897_wire;
      req(0) <= phi_stmt_1894_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1894_ack_0,
          idata => idata,
          odata => xx_xlcssa220_1894,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1894
    phi_stmt_1898: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1901_wire;
      req(0) <= phi_stmt_1898_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1898_ack_0,
          idata => idata,
          odata => xx_xlcssa219_1898,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1898
    phi_stmt_1902: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1905_wire;
      req(0) <= phi_stmt_1902_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1902_ack_0,
          idata => idata,
          odata => xx_xlcssa218_1902,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1902
    phi_stmt_1906: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1909_wire;
      req(0) <= phi_stmt_1906_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1906_ack_0,
          idata => idata,
          odata => xx_xlcssa217_1906,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1906
    phi_stmt_1910: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1913_wire;
      req(0) <= phi_stmt_1910_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1910_ack_0,
          idata => idata,
          odata => xx_xlcssa216_1910,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1910
    phi_stmt_1914: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1917_wire;
      req(0) <= phi_stmt_1914_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1914_ack_0,
          idata => idata,
          odata => xx_xlcssa215_1914,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1914
    phi_stmt_1918: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1921_wire;
      req(0) <= phi_stmt_1918_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1918_ack_0,
          idata => idata,
          odata => xx_xlcssa214_1918,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1918
    phi_stmt_1922: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1925_wire;
      req(0) <= phi_stmt_1922_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1922_ack_0,
          idata => idata,
          odata => xx_xlcssa213_1922,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1922
    phi_stmt_1926: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1929_wire;
      req(0) <= phi_stmt_1926_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1926_ack_0,
          idata => idata,
          odata => xx_xlcssa212_1926,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1926
    phi_stmt_1930: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1933_wire;
      req(0) <= phi_stmt_1930_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1930_ack_0,
          idata => idata,
          odata => xx_xlcssa211_1930,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1930
    phi_stmt_1934: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1937_wire;
      req(0) <= phi_stmt_1934_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1934_ack_0,
          idata => idata,
          odata => xx_xlcssa210_1934,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1934
    phi_stmt_1938: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1941_wire;
      req(0) <= phi_stmt_1938_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1938_ack_0,
          idata => idata,
          odata => xx_xlcssa209_1938,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1938
    phi_stmt_1942: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1945_wire;
      req(0) <= phi_stmt_1942_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1942_ack_0,
          idata => idata,
          odata => xx_xlcssa208_1942,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1942
    phi_stmt_1946: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1949_wire;
      req(0) <= phi_stmt_1946_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1946_ack_0,
          idata => idata,
          odata => xx_xlcssa207_1946,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1946
    phi_stmt_1950: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1953_wire;
      req(0) <= phi_stmt_1950_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1950_ack_0,
          idata => idata,
          odata => xx_xlcssa_1950,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1950
    phi_stmt_555: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_559_wire_constant & type_cast_561_wire;
      req <= phi_stmt_555_req_0 & phi_stmt_555_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_555_ack_0,
          idata => idata,
          odata => indvar60_555,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_555
    phi_stmt_589: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_593_wire_constant & type_cast_595_wire;
      req <= phi_stmt_589_req_0 & phi_stmt_589_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_589_ack_0,
          idata => idata,
          odata => indvar56_589,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_589
    phi_stmt_743: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_747_wire_constant & type_cast_749_wire;
      req <= phi_stmt_743_req_0 & phi_stmt_743_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_743_ack_0,
          idata => idata,
          odata => indvar_743,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_743
    phi_stmt_750: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_754_wire_constant & type_cast_756_wire;
      req <= phi_stmt_750_req_0 & phi_stmt_750_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_750_ack_0,
          idata => idata,
          odata => v33x_x018_750,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_750
    phi_stmt_757: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_761_wire_constant & type_cast_763_wire;
      req <= phi_stmt_757_req_0 & phi_stmt_757_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_757_ack_0,
          idata => idata,
          odata => v32x_x017_757,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_757
    phi_stmt_764: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_768_wire_constant & type_cast_770_wire;
      req <= phi_stmt_764_req_0 & phi_stmt_764_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_764_ack_0,
          idata => idata,
          odata => v31x_x016_764,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_764
    phi_stmt_771: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_775_wire_constant & type_cast_777_wire;
      req <= phi_stmt_771_req_0 & phi_stmt_771_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_771_ack_0,
          idata => idata,
          odata => v30x_x015_771,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_771
    phi_stmt_778: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_782_wire_constant & type_cast_784_wire;
      req <= phi_stmt_778_req_0 & phi_stmt_778_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_778_ack_0,
          idata => idata,
          odata => v23x_x014_778,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_778
    phi_stmt_785: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_789_wire_constant & type_cast_791_wire;
      req <= phi_stmt_785_req_0 & phi_stmt_785_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_785_ack_0,
          idata => idata,
          odata => v22x_x013_785,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_785
    phi_stmt_792: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_796_wire_constant & type_cast_798_wire;
      req <= phi_stmt_792_req_0 & phi_stmt_792_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_792_ack_0,
          idata => idata,
          odata => v21x_x012_792,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_792
    phi_stmt_799: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_803_wire_constant & type_cast_805_wire;
      req <= phi_stmt_799_req_0 & phi_stmt_799_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_799_ack_0,
          idata => idata,
          odata => v20x_x011_799,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_799
    phi_stmt_806: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_810_wire_constant & type_cast_812_wire;
      req <= phi_stmt_806_req_0 & phi_stmt_806_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_806_ack_0,
          idata => idata,
          odata => v13x_x010_806,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_806
    phi_stmt_813: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_817_wire_constant & type_cast_819_wire;
      req <= phi_stmt_813_req_0 & phi_stmt_813_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_813_ack_0,
          idata => idata,
          odata => v00x_x09_813,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_813
    phi_stmt_820: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_824_wire_constant & type_cast_826_wire;
      req <= phi_stmt_820_req_0 & phi_stmt_820_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_820_ack_0,
          idata => idata,
          odata => v01x_x08_820,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_820
    phi_stmt_827: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_831_wire_constant & type_cast_833_wire;
      req <= phi_stmt_827_req_0 & phi_stmt_827_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_827_ack_0,
          idata => idata,
          odata => v02x_x07_827,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_827
    phi_stmt_834: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_838_wire_constant & type_cast_840_wire;
      req <= phi_stmt_834_req_0 & phi_stmt_834_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_834_ack_0,
          idata => idata,
          odata => v03x_x06_834,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_834
    phi_stmt_841: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_845_wire_constant & type_cast_847_wire;
      req <= phi_stmt_841_req_0 & phi_stmt_841_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_841_ack_0,
          idata => idata,
          odata => v10x_x05_841,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_841
    phi_stmt_848: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_852_wire_constant & type_cast_854_wire;
      req <= phi_stmt_848_req_0 & phi_stmt_848_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_848_ack_0,
          idata => idata,
          odata => v11x_x04_848,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_848
    phi_stmt_855: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_859_wire_constant & type_cast_861_wire;
      req <= phi_stmt_855_req_0 & phi_stmt_855_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_855_ack_0,
          idata => idata,
          odata => v12x_x03_855,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_855
    register_block_0 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1011_final_reg_req_0;
      addr_of_1011_final_reg_ack_0 <= ack; 
      addr_of_1011_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1010_root_address, dout => scevgep89_1012, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_1 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1023_final_reg_req_0;
      addr_of_1023_final_reg_ack_0 <= ack; 
      addr_of_1023_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1022_root_address, dout => scevgep80_1024, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_2 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1029_final_reg_req_0;
      addr_of_1029_final_reg_ack_0 <= ack; 
      addr_of_1029_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1028_root_address, dout => scevgep69_1030, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_3 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1035_final_reg_req_0;
      addr_of_1035_final_reg_ack_0 <= ack; 
      addr_of_1035_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1034_root_address, dout => scevgep97_1036, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_4 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1041_final_reg_req_0;
      addr_of_1041_final_reg_ack_0 <= ack; 
      addr_of_1041_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1040_root_address, dout => scevgep88_1042, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_5 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1047_final_reg_req_0;
      addr_of_1047_final_reg_ack_0 <= ack; 
      addr_of_1047_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1046_root_address, dout => scevgep79_1048, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_6 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1053_final_reg_req_0;
      addr_of_1053_final_reg_ack_0 <= ack; 
      addr_of_1053_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1052_root_address, dout => scevgep68_1054, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_7 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1059_final_reg_req_0;
      addr_of_1059_final_reg_ack_0 <= ack; 
      addr_of_1059_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1058_root_address, dout => scevgep96_1060, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_8 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1065_final_reg_req_0;
      addr_of_1065_final_reg_ack_0 <= ack; 
      addr_of_1065_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1064_root_address, dout => scevgep87_1066, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_9 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1071_final_reg_req_0;
      addr_of_1071_final_reg_ack_0 <= ack; 
      addr_of_1071_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1070_root_address, dout => scevgep78_1072, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_10 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1077_final_reg_req_0;
      addr_of_1077_final_reg_ack_0 <= ack; 
      addr_of_1077_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1076_root_address, dout => scevgep66_1078, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_11 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1083_final_reg_req_0;
      addr_of_1083_final_reg_ack_0 <= ack; 
      addr_of_1083_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1082_root_address, dout => scevgep94_1084, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_12 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1089_final_reg_req_0;
      addr_of_1089_final_reg_ack_0 <= ack; 
      addr_of_1089_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1088_root_address, dout => scevgep85_1090, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_13 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1095_final_reg_req_0;
      addr_of_1095_final_reg_ack_0 <= ack; 
      addr_of_1095_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1094_root_address, dout => scevgep76_1096, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_14 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1101_final_reg_req_0;
      addr_of_1101_final_reg_ack_0 <= ack; 
      addr_of_1101_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_1100_root_address, dout => scevgep_1102, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_15 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_607_final_reg_req_0;
      addr_of_607_final_reg_ack_0 <= ack; 
      addr_of_607_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_606_root_address, dout => scevgep134_608, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_16 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_619_final_reg_req_0;
      addr_of_619_final_reg_ack_0 <= ack; 
      addr_of_619_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_618_root_address, dout => scevgep146_620, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_17 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_631_final_reg_req_0;
      addr_of_631_final_reg_ack_0 <= ack; 
      addr_of_631_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_630_root_address, dout => scevgep142_632, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_18 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_637_final_reg_req_0;
      addr_of_637_final_reg_ack_0 <= ack; 
      addr_of_637_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_636_root_address, dout => scevgep129_638, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_19 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_643_final_reg_req_0;
      addr_of_643_final_reg_ack_0 <= ack; 
      addr_of_643_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_642_root_address, dout => scevgep143_644, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_20 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_649_final_reg_req_0;
      addr_of_649_final_reg_ack_0 <= ack; 
      addr_of_649_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_648_root_address, dout => scevgep139_650, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_21 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_661_final_reg_req_0;
      addr_of_661_final_reg_ack_0 <= ack; 
      addr_of_661_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_660_root_address, dout => scevgep135_662, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_22 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_667_final_reg_req_0;
      addr_of_667_final_reg_ack_0 <= ack; 
      addr_of_667_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_666_root_address, dout => scevgep131_668, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_23 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_673_final_reg_req_0;
      addr_of_673_final_reg_ack_0 <= ack; 
      addr_of_673_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_672_root_address, dout => scevgep144_674, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_24 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_679_final_reg_req_0;
      addr_of_679_final_reg_ack_0 <= ack; 
      addr_of_679_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_678_root_address, dout => scevgep140_680, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_25 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_685_final_reg_req_0;
      addr_of_685_final_reg_ack_0 <= ack; 
      addr_of_685_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_684_root_address, dout => scevgep136_686, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_26 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_691_final_reg_req_0;
      addr_of_691_final_reg_ack_0 <= ack; 
      addr_of_691_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_690_root_address, dout => scevgep133_692, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_27 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_697_final_reg_req_0;
      addr_of_697_final_reg_ack_0 <= ack; 
      addr_of_697_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_696_root_address, dout => scevgep145_698, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_28 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_703_final_reg_req_0;
      addr_of_703_final_reg_ack_0 <= ack; 
      addr_of_703_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_702_root_address, dout => scevgep141_704, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_29 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_709_final_reg_req_0;
      addr_of_709_final_reg_ack_0 <= ack; 
      addr_of_709_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_708_root_address, dout => scevgep137_710, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_30 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_715_final_reg_req_0;
      addr_of_715_final_reg_ack_0 <= ack; 
      addr_of_715_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_714_root_address, dout => scevgep138_716, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_31 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_873_final_reg_req_0;
      addr_of_873_final_reg_ack_0 <= ack; 
      addr_of_873_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_872_root_address, dout => scevgep74_874, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_32 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_885_final_reg_req_0;
      addr_of_885_final_reg_ack_0 <= ack; 
      addr_of_885_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_884_root_address, dout => scevgep101_886, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_33 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_897_final_reg_req_0;
      addr_of_897_final_reg_ack_0 <= ack; 
      addr_of_897_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_896_root_address, dout => scevgep92_898, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_34 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_903_final_reg_req_0;
      addr_of_903_final_reg_ack_0 <= ack; 
      addr_of_903_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_902_root_address, dout => scevgep64_904, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_35 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_909_final_reg_req_0;
      addr_of_909_final_reg_ack_0 <= ack; 
      addr_of_909_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_908_root_address, dout => scevgep95_910, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_36 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_915_final_reg_req_0;
      addr_of_915_final_reg_ack_0 <= ack; 
      addr_of_915_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_914_root_address, dout => scevgep86_916, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_37 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_927_final_reg_req_0;
      addr_of_927_final_reg_ack_0 <= ack; 
      addr_of_927_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_926_root_address, dout => scevgep77_928, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_38 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_933_final_reg_req_0;
      addr_of_933_final_reg_ack_0 <= ack; 
      addr_of_933_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_932_root_address, dout => scevgep71_934, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_39 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_939_final_reg_req_0;
      addr_of_939_final_reg_ack_0 <= ack; 
      addr_of_939_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_938_root_address, dout => scevgep99_940, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_40 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_945_final_reg_req_0;
      addr_of_945_final_reg_ack_0 <= ack; 
      addr_of_945_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_944_root_address, dout => scevgep90_946, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_41 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_951_final_reg_req_0;
      addr_of_951_final_reg_ack_0 <= ack; 
      addr_of_951_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_950_root_address, dout => scevgep81_952, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_42 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_957_final_reg_req_0;
      addr_of_957_final_reg_ack_0 <= ack; 
      addr_of_957_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_956_root_address, dout => scevgep73_958, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_43 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_963_final_reg_req_0;
      addr_of_963_final_reg_ack_0 <= ack; 
      addr_of_963_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_962_root_address, dout => scevgep100_964, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_44 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_969_final_reg_req_0;
      addr_of_969_final_reg_ack_0 <= ack; 
      addr_of_969_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_968_root_address, dout => scevgep91_970, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_45 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_975_final_reg_req_0;
      addr_of_975_final_reg_ack_0 <= ack; 
      addr_of_975_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_974_root_address, dout => scevgep82_976, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_46 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_981_final_reg_req_0;
      addr_of_981_final_reg_ack_0 <= ack; 
      addr_of_981_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_980_root_address, dout => scevgep83_982, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_47 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_999_final_reg_req_0;
      addr_of_999_final_reg_ack_0 <= ack; 
      addr_of_999_final_reg: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 32) 
        port map( din => array_obj_ref_998_root_address, dout => scevgep98_1000, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_48 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1010_index_0_resize_req_0;
      array_obj_ref_1010_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1010_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp270_1006, dout => simple_obj_ref_1008_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_49 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1010_index_1_resize_req_0;
      array_obj_ref_1010_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1010_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp268_722, dout => simple_obj_ref_1009_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_50 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1010_offset_inst_req_0;
      array_obj_ref_1010_offset_inst_ack_0 <= ack; 
      array_obj_ref_1010_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1010_index_partial_sum_1, dout => array_obj_ref_1010_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_51 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1022_index_0_resize_req_0;
      array_obj_ref_1022_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1022_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp272_1018, dout => simple_obj_ref_1020_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_52 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1022_index_1_resize_req_0;
      array_obj_ref_1022_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1022_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp268_722, dout => simple_obj_ref_1021_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_53 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1022_offset_inst_req_0;
      array_obj_ref_1022_offset_inst_ack_0 <= ack; 
      array_obj_ref_1022_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1022_index_partial_sum_1, dout => array_obj_ref_1022_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_54 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1028_index_0_resize_req_0;
      array_obj_ref_1028_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1028_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp266_988, dout => simple_obj_ref_1026_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_55 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1028_index_1_resize_req_0;
      array_obj_ref_1028_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1028_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp268_722, dout => simple_obj_ref_1027_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_56 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1028_offset_inst_req_0;
      array_obj_ref_1028_offset_inst_ack_0 <= ack; 
      array_obj_ref_1028_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1028_index_partial_sum_1, dout => array_obj_ref_1028_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_57 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1034_index_0_resize_req_0;
      array_obj_ref_1034_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1034_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp267_994, dout => simple_obj_ref_1032_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_58 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1034_index_1_resize_req_0;
      array_obj_ref_1034_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1034_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp275_728, dout => simple_obj_ref_1033_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_59 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1034_offset_inst_req_0;
      array_obj_ref_1034_offset_inst_ack_0 <= ack; 
      array_obj_ref_1034_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1034_index_partial_sum_1, dout => array_obj_ref_1034_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_60 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1040_index_0_resize_req_0;
      array_obj_ref_1040_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1040_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp270_1006, dout => simple_obj_ref_1038_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_61 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1040_index_1_resize_req_0;
      array_obj_ref_1040_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1040_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp275_728, dout => simple_obj_ref_1039_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_62 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1040_offset_inst_req_0;
      array_obj_ref_1040_offset_inst_ack_0 <= ack; 
      array_obj_ref_1040_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1040_index_partial_sum_1, dout => array_obj_ref_1040_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_63 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1046_index_0_resize_req_0;
      array_obj_ref_1046_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1046_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp272_1018, dout => simple_obj_ref_1044_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_64 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1046_index_1_resize_req_0;
      array_obj_ref_1046_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1046_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp275_728, dout => simple_obj_ref_1045_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_65 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1046_offset_inst_req_0;
      array_obj_ref_1046_offset_inst_ack_0 <= ack; 
      array_obj_ref_1046_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1046_index_partial_sum_1, dout => array_obj_ref_1046_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_66 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1052_index_0_resize_req_0;
      array_obj_ref_1052_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1052_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp266_988, dout => simple_obj_ref_1050_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_67 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1052_index_1_resize_req_0;
      array_obj_ref_1052_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1052_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp275_728, dout => simple_obj_ref_1051_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_68 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1052_offset_inst_req_0;
      array_obj_ref_1052_offset_inst_ack_0 <= ack; 
      array_obj_ref_1052_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1052_index_partial_sum_1, dout => array_obj_ref_1052_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_69 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1058_index_0_resize_req_0;
      array_obj_ref_1058_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1058_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp267_994, dout => simple_obj_ref_1056_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_70 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1058_index_1_resize_req_0;
      array_obj_ref_1058_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1058_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp280_734, dout => simple_obj_ref_1057_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_71 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1058_offset_inst_req_0;
      array_obj_ref_1058_offset_inst_ack_0 <= ack; 
      array_obj_ref_1058_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1058_index_partial_sum_1, dout => array_obj_ref_1058_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_72 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1064_index_0_resize_req_0;
      array_obj_ref_1064_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1064_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp270_1006, dout => simple_obj_ref_1062_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_73 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1064_index_1_resize_req_0;
      array_obj_ref_1064_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1064_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp280_734, dout => simple_obj_ref_1063_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_74 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1064_offset_inst_req_0;
      array_obj_ref_1064_offset_inst_ack_0 <= ack; 
      array_obj_ref_1064_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1064_index_partial_sum_1, dout => array_obj_ref_1064_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_75 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1070_index_0_resize_req_0;
      array_obj_ref_1070_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1070_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp272_1018, dout => simple_obj_ref_1068_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_76 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1070_index_1_resize_req_0;
      array_obj_ref_1070_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1070_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp280_734, dout => simple_obj_ref_1069_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_77 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1070_offset_inst_req_0;
      array_obj_ref_1070_offset_inst_ack_0 <= ack; 
      array_obj_ref_1070_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1070_index_partial_sum_1, dout => array_obj_ref_1070_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_78 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1076_index_0_resize_req_0;
      array_obj_ref_1076_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1076_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp266_988, dout => simple_obj_ref_1074_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_79 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1076_index_1_resize_req_0;
      array_obj_ref_1076_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1076_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp280_734, dout => simple_obj_ref_1075_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_80 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1076_offset_inst_req_0;
      array_obj_ref_1076_offset_inst_ack_0 <= ack; 
      array_obj_ref_1076_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1076_index_partial_sum_1, dout => array_obj_ref_1076_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_81 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1082_index_0_resize_req_0;
      array_obj_ref_1082_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1082_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp267_994, dout => simple_obj_ref_1080_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_82 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1082_index_1_resize_req_0;
      array_obj_ref_1082_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1082_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp285_740, dout => simple_obj_ref_1081_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_83 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1082_offset_inst_req_0;
      array_obj_ref_1082_offset_inst_ack_0 <= ack; 
      array_obj_ref_1082_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1082_index_partial_sum_1, dout => array_obj_ref_1082_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_84 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1088_index_0_resize_req_0;
      array_obj_ref_1088_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1088_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp270_1006, dout => simple_obj_ref_1086_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_85 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1088_index_1_resize_req_0;
      array_obj_ref_1088_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1088_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp285_740, dout => simple_obj_ref_1087_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_86 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1088_offset_inst_req_0;
      array_obj_ref_1088_offset_inst_ack_0 <= ack; 
      array_obj_ref_1088_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1088_index_partial_sum_1, dout => array_obj_ref_1088_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_87 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1094_index_0_resize_req_0;
      array_obj_ref_1094_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1094_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp272_1018, dout => simple_obj_ref_1092_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_88 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1094_index_1_resize_req_0;
      array_obj_ref_1094_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1094_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp285_740, dout => simple_obj_ref_1093_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_89 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1094_offset_inst_req_0;
      array_obj_ref_1094_offset_inst_ack_0 <= ack; 
      array_obj_ref_1094_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1094_index_partial_sum_1, dout => array_obj_ref_1094_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_90 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1100_index_0_resize_req_0;
      array_obj_ref_1100_index_0_resize_ack_0 <= ack; 
      array_obj_ref_1100_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp266_988, dout => simple_obj_ref_1098_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_91 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1100_index_1_resize_req_0;
      array_obj_ref_1100_index_1_resize_ack_0 <= ack; 
      array_obj_ref_1100_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp285_740, dout => simple_obj_ref_1099_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_92 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_1100_offset_inst_req_0;
      array_obj_ref_1100_offset_inst_ack_0 <= ack; 
      array_obj_ref_1100_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_1100_index_partial_sum_1, dout => array_obj_ref_1100_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_93 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_606_index_0_resize_req_0;
      array_obj_ref_606_index_0_resize_ack_0 <= ack; 
      array_obj_ref_606_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_604_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_94 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_606_index_1_resize_req_0;
      array_obj_ref_606_index_1_resize_ack_0 <= ack; 
      array_obj_ref_606_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp312_602, dout => simple_obj_ref_605_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_95 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_606_offset_inst_req_0;
      array_obj_ref_606_offset_inst_ack_0 <= ack; 
      array_obj_ref_606_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_606_index_partial_sum_1, dout => array_obj_ref_606_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_96 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_618_index_0_resize_req_0;
      array_obj_ref_618_index_0_resize_ack_0 <= ack; 
      array_obj_ref_618_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_616_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_97 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_618_index_1_resize_req_0;
      array_obj_ref_618_index_1_resize_ack_0 <= ack; 
      array_obj_ref_618_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp314_614, dout => simple_obj_ref_617_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_98 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_618_offset_inst_req_0;
      array_obj_ref_618_offset_inst_ack_0 <= ack; 
      array_obj_ref_618_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_618_index_partial_sum_1, dout => array_obj_ref_618_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_99 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_630_index_0_resize_req_0;
      array_obj_ref_630_index_0_resize_ack_0 <= ack; 
      array_obj_ref_630_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_628_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_100 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_630_index_1_resize_req_0;
      array_obj_ref_630_index_1_resize_ack_0 <= ack; 
      array_obj_ref_630_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp316_626, dout => simple_obj_ref_629_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_101 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_630_offset_inst_req_0;
      array_obj_ref_630_offset_inst_ack_0 <= ack; 
      array_obj_ref_630_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_630_index_partial_sum_1, dout => array_obj_ref_630_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_102 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_636_index_0_resize_req_0;
      array_obj_ref_636_index_0_resize_ack_0 <= ack; 
      array_obj_ref_636_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_634_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_103 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_636_index_1_resize_req_0;
      array_obj_ref_636_index_1_resize_ack_0 <= ack; 
      array_obj_ref_636_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp312_602, dout => simple_obj_ref_635_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_104 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_636_offset_inst_req_0;
      array_obj_ref_636_offset_inst_ack_0 <= ack; 
      array_obj_ref_636_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_636_index_partial_sum_1, dout => array_obj_ref_636_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_105 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_642_index_0_resize_req_0;
      array_obj_ref_642_index_0_resize_ack_0 <= ack; 
      array_obj_ref_642_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_640_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_106 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_642_index_1_resize_req_0;
      array_obj_ref_642_index_1_resize_ack_0 <= ack; 
      array_obj_ref_642_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp314_614, dout => simple_obj_ref_641_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_107 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_642_offset_inst_req_0;
      array_obj_ref_642_offset_inst_ack_0 <= ack; 
      array_obj_ref_642_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_642_index_partial_sum_1, dout => array_obj_ref_642_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_108 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_648_index_0_resize_req_0;
      array_obj_ref_648_index_0_resize_ack_0 <= ack; 
      array_obj_ref_648_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_646_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_109 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_648_index_1_resize_req_0;
      array_obj_ref_648_index_1_resize_ack_0 <= ack; 
      array_obj_ref_648_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp316_626, dout => simple_obj_ref_647_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_110 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_648_offset_inst_req_0;
      array_obj_ref_648_offset_inst_ack_0 <= ack; 
      array_obj_ref_648_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_648_index_partial_sum_1, dout => array_obj_ref_648_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_111 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_660_index_0_resize_req_0;
      array_obj_ref_660_index_0_resize_ack_0 <= ack; 
      array_obj_ref_660_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_658_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_112 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_660_index_1_resize_req_0;
      array_obj_ref_660_index_1_resize_ack_0 <= ack; 
      array_obj_ref_660_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp322_656, dout => simple_obj_ref_659_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_113 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_660_offset_inst_req_0;
      array_obj_ref_660_offset_inst_ack_0 <= ack; 
      array_obj_ref_660_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_660_index_partial_sum_1, dout => array_obj_ref_660_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_114 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_666_index_0_resize_req_0;
      array_obj_ref_666_index_0_resize_ack_0 <= ack; 
      array_obj_ref_666_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_664_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_115 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_666_index_1_resize_req_0;
      array_obj_ref_666_index_1_resize_ack_0 <= ack; 
      array_obj_ref_666_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp312_602, dout => simple_obj_ref_665_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_116 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_666_offset_inst_req_0;
      array_obj_ref_666_offset_inst_ack_0 <= ack; 
      array_obj_ref_666_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_666_index_partial_sum_1, dout => array_obj_ref_666_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_117 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_672_index_0_resize_req_0;
      array_obj_ref_672_index_0_resize_ack_0 <= ack; 
      array_obj_ref_672_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_670_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_118 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_672_index_1_resize_req_0;
      array_obj_ref_672_index_1_resize_ack_0 <= ack; 
      array_obj_ref_672_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp314_614, dout => simple_obj_ref_671_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_119 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_672_offset_inst_req_0;
      array_obj_ref_672_offset_inst_ack_0 <= ack; 
      array_obj_ref_672_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_672_index_partial_sum_1, dout => array_obj_ref_672_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_120 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_678_index_0_resize_req_0;
      array_obj_ref_678_index_0_resize_ack_0 <= ack; 
      array_obj_ref_678_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_676_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_121 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_678_index_1_resize_req_0;
      array_obj_ref_678_index_1_resize_ack_0 <= ack; 
      array_obj_ref_678_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp316_626, dout => simple_obj_ref_677_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_122 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_678_offset_inst_req_0;
      array_obj_ref_678_offset_inst_ack_0 <= ack; 
      array_obj_ref_678_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_678_index_partial_sum_1, dout => array_obj_ref_678_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_123 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_684_index_0_resize_req_0;
      array_obj_ref_684_index_0_resize_ack_0 <= ack; 
      array_obj_ref_684_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_682_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_124 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_684_index_1_resize_req_0;
      array_obj_ref_684_index_1_resize_ack_0 <= ack; 
      array_obj_ref_684_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp322_656, dout => simple_obj_ref_683_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_125 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_684_offset_inst_req_0;
      array_obj_ref_684_offset_inst_ack_0 <= ack; 
      array_obj_ref_684_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_684_index_partial_sum_1, dout => array_obj_ref_684_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_126 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_690_index_0_resize_req_0;
      array_obj_ref_690_index_0_resize_ack_0 <= ack; 
      array_obj_ref_690_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_688_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_127 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_690_index_1_resize_req_0;
      array_obj_ref_690_index_1_resize_ack_0 <= ack; 
      array_obj_ref_690_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp312_602, dout => simple_obj_ref_689_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_128 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_690_offset_inst_req_0;
      array_obj_ref_690_offset_inst_ack_0 <= ack; 
      array_obj_ref_690_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_690_index_partial_sum_1, dout => array_obj_ref_690_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_129 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_696_index_0_resize_req_0;
      array_obj_ref_696_index_0_resize_ack_0 <= ack; 
      array_obj_ref_696_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_694_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_130 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_696_index_1_resize_req_0;
      array_obj_ref_696_index_1_resize_ack_0 <= ack; 
      array_obj_ref_696_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp314_614, dout => simple_obj_ref_695_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_131 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_696_offset_inst_req_0;
      array_obj_ref_696_offset_inst_ack_0 <= ack; 
      array_obj_ref_696_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_696_index_partial_sum_1, dout => array_obj_ref_696_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_132 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_702_index_0_resize_req_0;
      array_obj_ref_702_index_0_resize_ack_0 <= ack; 
      array_obj_ref_702_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_700_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_133 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_702_index_1_resize_req_0;
      array_obj_ref_702_index_1_resize_ack_0 <= ack; 
      array_obj_ref_702_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp316_626, dout => simple_obj_ref_701_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_134 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_702_offset_inst_req_0;
      array_obj_ref_702_offset_inst_ack_0 <= ack; 
      array_obj_ref_702_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_702_index_partial_sum_1, dout => array_obj_ref_702_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_135 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_708_index_0_resize_req_0;
      array_obj_ref_708_index_0_resize_ack_0 <= ack; 
      array_obj_ref_708_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_706_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_136 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_708_index_1_resize_req_0;
      array_obj_ref_708_index_1_resize_ack_0 <= ack; 
      array_obj_ref_708_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp322_656, dout => simple_obj_ref_707_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_137 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_708_offset_inst_req_0;
      array_obj_ref_708_offset_inst_ack_0 <= ack; 
      array_obj_ref_708_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_708_index_partial_sum_1, dout => array_obj_ref_708_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_138 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_714_index_0_resize_req_0;
      array_obj_ref_714_index_0_resize_ack_0 <= ack; 
      array_obj_ref_714_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_712_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_139 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_714_index_1_resize_req_0;
      array_obj_ref_714_index_1_resize_ack_0 <= ack; 
      array_obj_ref_714_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp322_656, dout => simple_obj_ref_713_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_140 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_714_offset_inst_req_0;
      array_obj_ref_714_offset_inst_ack_0 <= ack; 
      array_obj_ref_714_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_714_index_partial_sum_1, dout => array_obj_ref_714_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_141 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_872_index_0_resize_req_0;
      array_obj_ref_872_index_0_resize_ack_0 <= ack; 
      array_obj_ref_872_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_870_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_142 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_872_index_1_resize_req_0;
      array_obj_ref_872_index_1_resize_ack_0 <= ack; 
      array_obj_ref_872_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp335_868, dout => simple_obj_ref_871_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_143 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_872_offset_inst_req_0;
      array_obj_ref_872_offset_inst_ack_0 <= ack; 
      array_obj_ref_872_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_872_index_partial_sum_1, dout => array_obj_ref_872_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_144 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_884_index_0_resize_req_0;
      array_obj_ref_884_index_0_resize_ack_0 <= ack; 
      array_obj_ref_884_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_882_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_145 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_884_index_1_resize_req_0;
      array_obj_ref_884_index_1_resize_ack_0 <= ack; 
      array_obj_ref_884_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp337_880, dout => simple_obj_ref_883_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_146 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_884_offset_inst_req_0;
      array_obj_ref_884_offset_inst_ack_0 <= ack; 
      array_obj_ref_884_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_884_index_partial_sum_1, dout => array_obj_ref_884_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_147 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_896_index_0_resize_req_0;
      array_obj_ref_896_index_0_resize_ack_0 <= ack; 
      array_obj_ref_896_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_894_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_148 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_896_index_1_resize_req_0;
      array_obj_ref_896_index_1_resize_ack_0 <= ack; 
      array_obj_ref_896_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp339_892, dout => simple_obj_ref_895_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_149 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_896_offset_inst_req_0;
      array_obj_ref_896_offset_inst_ack_0 <= ack; 
      array_obj_ref_896_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_896_index_partial_sum_1, dout => array_obj_ref_896_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_150 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_902_index_0_resize_req_0;
      array_obj_ref_902_index_0_resize_ack_0 <= ack; 
      array_obj_ref_902_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_900_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_151 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_902_index_1_resize_req_0;
      array_obj_ref_902_index_1_resize_ack_0 <= ack; 
      array_obj_ref_902_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp335_868, dout => simple_obj_ref_901_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_152 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_902_offset_inst_req_0;
      array_obj_ref_902_offset_inst_ack_0 <= ack; 
      array_obj_ref_902_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_902_index_partial_sum_1, dout => array_obj_ref_902_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_153 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_908_index_0_resize_req_0;
      array_obj_ref_908_index_0_resize_ack_0 <= ack; 
      array_obj_ref_908_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_906_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_154 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_908_index_1_resize_req_0;
      array_obj_ref_908_index_1_resize_ack_0 <= ack; 
      array_obj_ref_908_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp337_880, dout => simple_obj_ref_907_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_155 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_908_offset_inst_req_0;
      array_obj_ref_908_offset_inst_ack_0 <= ack; 
      array_obj_ref_908_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_908_index_partial_sum_1, dout => array_obj_ref_908_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_156 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_914_index_0_resize_req_0;
      array_obj_ref_914_index_0_resize_ack_0 <= ack; 
      array_obj_ref_914_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_912_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_157 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_914_index_1_resize_req_0;
      array_obj_ref_914_index_1_resize_ack_0 <= ack; 
      array_obj_ref_914_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp339_892, dout => simple_obj_ref_913_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_158 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_914_offset_inst_req_0;
      array_obj_ref_914_offset_inst_ack_0 <= ack; 
      array_obj_ref_914_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_914_index_partial_sum_1, dout => array_obj_ref_914_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_159 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_926_index_0_resize_req_0;
      array_obj_ref_926_index_0_resize_ack_0 <= ack; 
      array_obj_ref_926_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp318_574, dout => simple_obj_ref_924_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_160 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_926_index_1_resize_req_0;
      array_obj_ref_926_index_1_resize_ack_0 <= ack; 
      array_obj_ref_926_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp344_922, dout => simple_obj_ref_925_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_161 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_926_offset_inst_req_0;
      array_obj_ref_926_offset_inst_ack_0 <= ack; 
      array_obj_ref_926_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_926_index_partial_sum_1, dout => array_obj_ref_926_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_162 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_932_index_0_resize_req_0;
      array_obj_ref_932_index_0_resize_ack_0 <= ack; 
      array_obj_ref_932_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_930_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_163 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_932_index_1_resize_req_0;
      array_obj_ref_932_index_1_resize_ack_0 <= ack; 
      array_obj_ref_932_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp335_868, dout => simple_obj_ref_931_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_164 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_932_offset_inst_req_0;
      array_obj_ref_932_offset_inst_ack_0 <= ack; 
      array_obj_ref_932_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_932_index_partial_sum_1, dout => array_obj_ref_932_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_165 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_938_index_0_resize_req_0;
      array_obj_ref_938_index_0_resize_ack_0 <= ack; 
      array_obj_ref_938_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_936_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_166 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_938_index_1_resize_req_0;
      array_obj_ref_938_index_1_resize_ack_0 <= ack; 
      array_obj_ref_938_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp337_880, dout => simple_obj_ref_937_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_167 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_938_offset_inst_req_0;
      array_obj_ref_938_offset_inst_ack_0 <= ack; 
      array_obj_ref_938_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_938_index_partial_sum_1, dout => array_obj_ref_938_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_168 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_944_index_0_resize_req_0;
      array_obj_ref_944_index_0_resize_ack_0 <= ack; 
      array_obj_ref_944_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_942_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_169 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_944_index_1_resize_req_0;
      array_obj_ref_944_index_1_resize_ack_0 <= ack; 
      array_obj_ref_944_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp339_892, dout => simple_obj_ref_943_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_170 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_944_offset_inst_req_0;
      array_obj_ref_944_offset_inst_ack_0 <= ack; 
      array_obj_ref_944_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_944_index_partial_sum_1, dout => array_obj_ref_944_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_171 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_950_index_0_resize_req_0;
      array_obj_ref_950_index_0_resize_ack_0 <= ack; 
      array_obj_ref_950_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp324_580, dout => simple_obj_ref_948_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_172 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_950_index_1_resize_req_0;
      array_obj_ref_950_index_1_resize_ack_0 <= ack; 
      array_obj_ref_950_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp344_922, dout => simple_obj_ref_949_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_173 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_950_offset_inst_req_0;
      array_obj_ref_950_offset_inst_ack_0 <= ack; 
      array_obj_ref_950_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_950_index_partial_sum_1, dout => array_obj_ref_950_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_174 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_956_index_0_resize_req_0;
      array_obj_ref_956_index_0_resize_ack_0 <= ack; 
      array_obj_ref_956_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_954_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_175 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_956_index_1_resize_req_0;
      array_obj_ref_956_index_1_resize_ack_0 <= ack; 
      array_obj_ref_956_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp335_868, dout => simple_obj_ref_955_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_176 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_956_offset_inst_req_0;
      array_obj_ref_956_offset_inst_ack_0 <= ack; 
      array_obj_ref_956_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_956_index_partial_sum_1, dout => array_obj_ref_956_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_177 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_962_index_0_resize_req_0;
      array_obj_ref_962_index_0_resize_ack_0 <= ack; 
      array_obj_ref_962_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_960_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_178 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_962_index_1_resize_req_0;
      array_obj_ref_962_index_1_resize_ack_0 <= ack; 
      array_obj_ref_962_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp337_880, dout => simple_obj_ref_961_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_179 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_962_offset_inst_req_0;
      array_obj_ref_962_offset_inst_ack_0 <= ack; 
      array_obj_ref_962_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_962_index_partial_sum_1, dout => array_obj_ref_962_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_180 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_968_index_0_resize_req_0;
      array_obj_ref_968_index_0_resize_ack_0 <= ack; 
      array_obj_ref_968_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_966_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_181 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_968_index_1_resize_req_0;
      array_obj_ref_968_index_1_resize_ack_0 <= ack; 
      array_obj_ref_968_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp339_892, dout => simple_obj_ref_967_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_182 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_968_offset_inst_req_0;
      array_obj_ref_968_offset_inst_ack_0 <= ack; 
      array_obj_ref_968_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_968_index_partial_sum_1, dout => array_obj_ref_968_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_183 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_974_index_0_resize_req_0;
      array_obj_ref_974_index_0_resize_ack_0 <= ack; 
      array_obj_ref_974_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp329_586, dout => simple_obj_ref_972_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_184 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_974_index_1_resize_req_0;
      array_obj_ref_974_index_1_resize_ack_0 <= ack; 
      array_obj_ref_974_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp344_922, dout => simple_obj_ref_973_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_185 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_974_offset_inst_req_0;
      array_obj_ref_974_offset_inst_ack_0 <= ack; 
      array_obj_ref_974_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_974_index_partial_sum_1, dout => array_obj_ref_974_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_186 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_980_index_0_resize_req_0;
      array_obj_ref_980_index_0_resize_ack_0 <= ack; 
      array_obj_ref_980_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp311_568, dout => simple_obj_ref_978_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_187 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_980_index_1_resize_req_0;
      array_obj_ref_980_index_1_resize_ack_0 <= ack; 
      array_obj_ref_980_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp344_922, dout => simple_obj_ref_979_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_188 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_980_offset_inst_req_0;
      array_obj_ref_980_offset_inst_ack_0 <= ack; 
      array_obj_ref_980_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_980_index_partial_sum_1, dout => array_obj_ref_980_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_189 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_998_index_0_resize_req_0;
      array_obj_ref_998_index_0_resize_ack_0 <= ack; 
      array_obj_ref_998_index_0_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp267_994, dout => simple_obj_ref_996_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_190 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_998_index_1_resize_req_0;
      array_obj_ref_998_index_1_resize_ack_0 <= ack; 
      array_obj_ref_998_index_1_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => tmp268_722, dout => simple_obj_ref_997_resized, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_191 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= array_obj_ref_998_offset_inst_req_0;
      array_obj_ref_998_offset_inst_ack_0 <= ack; 
      array_obj_ref_998_offset_inst: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => array_obj_ref_998_index_partial_sum_1, dout => array_obj_ref_998_final_offset, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_192 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1105_addr_0_req_0;
      ptr_deref_1105_addr_0_ack_0 <= ack; 
      ptr_deref_1105_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1105_root_address, dout => ptr_deref_1105_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_193 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1105_base_resize_req_0;
      ptr_deref_1105_base_resize_ack_0 <= ack; 
      ptr_deref_1105_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep74_874, dout => ptr_deref_1105_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_194 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1109_addr_0_req_0;
      ptr_deref_1109_addr_0_ack_0 <= ack; 
      ptr_deref_1109_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1109_root_address, dout => ptr_deref_1109_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_195 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1109_base_resize_req_0;
      ptr_deref_1109_base_resize_ack_0 <= ack; 
      ptr_deref_1109_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep69_1030, dout => ptr_deref_1109_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_196 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1113_addr_0_req_0;
      ptr_deref_1113_addr_0_ack_0 <= ack; 
      ptr_deref_1113_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1113_root_address, dout => ptr_deref_1113_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_197 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1113_base_resize_req_0;
      ptr_deref_1113_base_resize_ack_0 <= ack; 
      ptr_deref_1113_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep83_982, dout => ptr_deref_1113_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_198 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1117_addr_0_req_0;
      ptr_deref_1117_addr_0_ack_0 <= ack; 
      ptr_deref_1117_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1117_root_address, dout => ptr_deref_1117_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_199 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1117_base_resize_req_0;
      ptr_deref_1117_base_resize_ack_0 <= ack; 
      ptr_deref_1117_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep80_1024, dout => ptr_deref_1117_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_200 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1121_addr_0_req_0;
      ptr_deref_1121_addr_0_ack_0 <= ack; 
      ptr_deref_1121_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1121_root_address, dout => ptr_deref_1121_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_201 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1121_base_resize_req_0;
      ptr_deref_1121_base_resize_ack_0 <= ack; 
      ptr_deref_1121_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep92_898, dout => ptr_deref_1121_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_202 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1125_addr_0_req_0;
      ptr_deref_1125_addr_0_ack_0 <= ack; 
      ptr_deref_1125_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1125_root_address, dout => ptr_deref_1125_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_203 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1125_base_resize_req_0;
      ptr_deref_1125_base_resize_ack_0 <= ack; 
      ptr_deref_1125_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep89_1012, dout => ptr_deref_1125_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_204 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1129_addr_0_req_0;
      ptr_deref_1129_addr_0_ack_0 <= ack; 
      ptr_deref_1129_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1129_root_address, dout => ptr_deref_1129_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_205 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1129_base_resize_req_0;
      ptr_deref_1129_base_resize_ack_0 <= ack; 
      ptr_deref_1129_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep101_886, dout => ptr_deref_1129_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_206 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1133_addr_0_req_0;
      ptr_deref_1133_addr_0_ack_0 <= ack; 
      ptr_deref_1133_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1133_root_address, dout => ptr_deref_1133_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_207 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1133_base_resize_req_0;
      ptr_deref_1133_base_resize_ack_0 <= ack; 
      ptr_deref_1133_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep98_1000, dout => ptr_deref_1133_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_208 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1177_addr_0_req_0;
      ptr_deref_1177_addr_0_ack_0 <= ack; 
      ptr_deref_1177_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1177_root_address, dout => ptr_deref_1177_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_209 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1177_base_resize_req_0;
      ptr_deref_1177_base_resize_ack_0 <= ack; 
      ptr_deref_1177_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep68_1054, dout => ptr_deref_1177_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_210 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1181_addr_0_req_0;
      ptr_deref_1181_addr_0_ack_0 <= ack; 
      ptr_deref_1181_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1181_root_address, dout => ptr_deref_1181_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_211 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1181_base_resize_req_0;
      ptr_deref_1181_base_resize_ack_0 <= ack; 
      ptr_deref_1181_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep79_1048, dout => ptr_deref_1181_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_212 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1185_addr_0_req_0;
      ptr_deref_1185_addr_0_ack_0 <= ack; 
      ptr_deref_1185_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1185_root_address, dout => ptr_deref_1185_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_213 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1185_base_resize_req_0;
      ptr_deref_1185_base_resize_ack_0 <= ack; 
      ptr_deref_1185_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep88_1042, dout => ptr_deref_1185_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_214 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1189_addr_0_req_0;
      ptr_deref_1189_addr_0_ack_0 <= ack; 
      ptr_deref_1189_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1189_root_address, dout => ptr_deref_1189_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_215 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1189_base_resize_req_0;
      ptr_deref_1189_base_resize_ack_0 <= ack; 
      ptr_deref_1189_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep97_1036, dout => ptr_deref_1189_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_216 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1233_addr_0_req_0;
      ptr_deref_1233_addr_0_ack_0 <= ack; 
      ptr_deref_1233_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1233_root_address, dout => ptr_deref_1233_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_217 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1233_base_resize_req_0;
      ptr_deref_1233_base_resize_ack_0 <= ack; 
      ptr_deref_1233_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep66_1078, dout => ptr_deref_1233_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_218 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1237_addr_0_req_0;
      ptr_deref_1237_addr_0_ack_0 <= ack; 
      ptr_deref_1237_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1237_root_address, dout => ptr_deref_1237_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_219 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1237_base_resize_req_0;
      ptr_deref_1237_base_resize_ack_0 <= ack; 
      ptr_deref_1237_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep78_1072, dout => ptr_deref_1237_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_220 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1241_addr_0_req_0;
      ptr_deref_1241_addr_0_ack_0 <= ack; 
      ptr_deref_1241_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1241_root_address, dout => ptr_deref_1241_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_221 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1241_base_resize_req_0;
      ptr_deref_1241_base_resize_ack_0 <= ack; 
      ptr_deref_1241_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep87_1066, dout => ptr_deref_1241_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_222 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1245_addr_0_req_0;
      ptr_deref_1245_addr_0_ack_0 <= ack; 
      ptr_deref_1245_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1245_root_address, dout => ptr_deref_1245_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_223 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1245_base_resize_req_0;
      ptr_deref_1245_base_resize_ack_0 <= ack; 
      ptr_deref_1245_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep96_1060, dout => ptr_deref_1245_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_224 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1289_addr_0_req_0;
      ptr_deref_1289_addr_0_ack_0 <= ack; 
      ptr_deref_1289_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1289_root_address, dout => ptr_deref_1289_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_225 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1289_base_resize_req_0;
      ptr_deref_1289_base_resize_ack_0 <= ack; 
      ptr_deref_1289_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep_1102, dout => ptr_deref_1289_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_226 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1293_addr_0_req_0;
      ptr_deref_1293_addr_0_ack_0 <= ack; 
      ptr_deref_1293_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1293_root_address, dout => ptr_deref_1293_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_227 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1293_base_resize_req_0;
      ptr_deref_1293_base_resize_ack_0 <= ack; 
      ptr_deref_1293_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep76_1096, dout => ptr_deref_1293_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_228 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1297_addr_0_req_0;
      ptr_deref_1297_addr_0_ack_0 <= ack; 
      ptr_deref_1297_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1297_root_address, dout => ptr_deref_1297_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_229 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1297_base_resize_req_0;
      ptr_deref_1297_base_resize_ack_0 <= ack; 
      ptr_deref_1297_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep85_1090, dout => ptr_deref_1297_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_230 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1301_addr_0_req_0;
      ptr_deref_1301_addr_0_ack_0 <= ack; 
      ptr_deref_1301_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1301_root_address, dout => ptr_deref_1301_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_231 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1301_base_resize_req_0;
      ptr_deref_1301_base_resize_ack_0 <= ack; 
      ptr_deref_1301_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep94_1084, dout => ptr_deref_1301_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_232 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1345_addr_0_req_0;
      ptr_deref_1345_addr_0_ack_0 <= ack; 
      ptr_deref_1345_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1345_root_address, dout => ptr_deref_1345_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_233 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1345_base_resize_req_0;
      ptr_deref_1345_base_resize_ack_0 <= ack; 
      ptr_deref_1345_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep73_958, dout => ptr_deref_1345_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_234 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1349_addr_0_req_0;
      ptr_deref_1349_addr_0_ack_0 <= ack; 
      ptr_deref_1349_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1349_root_address, dout => ptr_deref_1349_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_235 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1349_base_resize_req_0;
      ptr_deref_1349_base_resize_ack_0 <= ack; 
      ptr_deref_1349_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep82_976, dout => ptr_deref_1349_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_236 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1353_addr_0_req_0;
      ptr_deref_1353_addr_0_ack_0 <= ack; 
      ptr_deref_1353_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1353_root_address, dout => ptr_deref_1353_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_237 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1353_base_resize_req_0;
      ptr_deref_1353_base_resize_ack_0 <= ack; 
      ptr_deref_1353_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep91_970, dout => ptr_deref_1353_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_238 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1357_addr_0_req_0;
      ptr_deref_1357_addr_0_ack_0 <= ack; 
      ptr_deref_1357_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1357_root_address, dout => ptr_deref_1357_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_239 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1357_base_resize_req_0;
      ptr_deref_1357_base_resize_ack_0 <= ack; 
      ptr_deref_1357_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep100_964, dout => ptr_deref_1357_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_240 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1521_addr_0_req_0;
      ptr_deref_1521_addr_0_ack_0 <= ack; 
      ptr_deref_1521_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1521_root_address, dout => ptr_deref_1521_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_241 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1521_base_resize_req_0;
      ptr_deref_1521_base_resize_ack_0 <= ack; 
      ptr_deref_1521_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep71_934, dout => ptr_deref_1521_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_242 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1525_addr_0_req_0;
      ptr_deref_1525_addr_0_ack_0 <= ack; 
      ptr_deref_1525_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1525_root_address, dout => ptr_deref_1525_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_243 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1525_base_resize_req_0;
      ptr_deref_1525_base_resize_ack_0 <= ack; 
      ptr_deref_1525_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep81_952, dout => ptr_deref_1525_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_244 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1529_addr_0_req_0;
      ptr_deref_1529_addr_0_ack_0 <= ack; 
      ptr_deref_1529_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1529_root_address, dout => ptr_deref_1529_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_245 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1529_base_resize_req_0;
      ptr_deref_1529_base_resize_ack_0 <= ack; 
      ptr_deref_1529_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep90_946, dout => ptr_deref_1529_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_246 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1533_addr_0_req_0;
      ptr_deref_1533_addr_0_ack_0 <= ack; 
      ptr_deref_1533_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1533_root_address, dout => ptr_deref_1533_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_247 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1533_base_resize_req_0;
      ptr_deref_1533_base_resize_ack_0 <= ack; 
      ptr_deref_1533_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep99_940, dout => ptr_deref_1533_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_248 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1697_addr_0_req_0;
      ptr_deref_1697_addr_0_ack_0 <= ack; 
      ptr_deref_1697_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1697_root_address, dout => ptr_deref_1697_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_249 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1697_base_resize_req_0;
      ptr_deref_1697_base_resize_ack_0 <= ack; 
      ptr_deref_1697_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep64_904, dout => ptr_deref_1697_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_250 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1701_addr_0_req_0;
      ptr_deref_1701_addr_0_ack_0 <= ack; 
      ptr_deref_1701_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1701_root_address, dout => ptr_deref_1701_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_251 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1701_base_resize_req_0;
      ptr_deref_1701_base_resize_ack_0 <= ack; 
      ptr_deref_1701_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep77_928, dout => ptr_deref_1701_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_252 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1705_addr_0_req_0;
      ptr_deref_1705_addr_0_ack_0 <= ack; 
      ptr_deref_1705_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1705_root_address, dout => ptr_deref_1705_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_253 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1705_base_resize_req_0;
      ptr_deref_1705_base_resize_ack_0 <= ack; 
      ptr_deref_1705_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep86_916, dout => ptr_deref_1705_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_254 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1709_addr_0_req_0;
      ptr_deref_1709_addr_0_ack_0 <= ack; 
      ptr_deref_1709_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1709_root_address, dout => ptr_deref_1709_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_255 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1709_base_resize_req_0;
      ptr_deref_1709_base_resize_ack_0 <= ack; 
      ptr_deref_1709_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep95_910, dout => ptr_deref_1709_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_256 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1956_addr_0_req_0;
      ptr_deref_1956_addr_0_ack_0 <= ack; 
      ptr_deref_1956_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1956_root_address, dout => ptr_deref_1956_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_257 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1956_base_resize_req_0;
      ptr_deref_1956_base_resize_ack_0 <= ack; 
      ptr_deref_1956_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep134_608, dout => ptr_deref_1956_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_258 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1960_addr_0_req_0;
      ptr_deref_1960_addr_0_ack_0 <= ack; 
      ptr_deref_1960_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1960_root_address, dout => ptr_deref_1960_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_259 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1960_base_resize_req_0;
      ptr_deref_1960_base_resize_ack_0 <= ack; 
      ptr_deref_1960_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep138_716, dout => ptr_deref_1960_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_260 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1964_addr_0_req_0;
      ptr_deref_1964_addr_0_ack_0 <= ack; 
      ptr_deref_1964_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1964_root_address, dout => ptr_deref_1964_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_261 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1964_base_resize_req_0;
      ptr_deref_1964_base_resize_ack_0 <= ack; 
      ptr_deref_1964_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep142_632, dout => ptr_deref_1964_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_262 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1968_addr_0_req_0;
      ptr_deref_1968_addr_0_ack_0 <= ack; 
      ptr_deref_1968_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1968_root_address, dout => ptr_deref_1968_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_263 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1968_base_resize_req_0;
      ptr_deref_1968_base_resize_ack_0 <= ack; 
      ptr_deref_1968_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep146_620, dout => ptr_deref_1968_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_264 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1972_addr_0_req_0;
      ptr_deref_1972_addr_0_ack_0 <= ack; 
      ptr_deref_1972_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1972_root_address, dout => ptr_deref_1972_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_265 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1972_base_resize_req_0;
      ptr_deref_1972_base_resize_ack_0 <= ack; 
      ptr_deref_1972_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep133_692, dout => ptr_deref_1972_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_266 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1976_addr_0_req_0;
      ptr_deref_1976_addr_0_ack_0 <= ack; 
      ptr_deref_1976_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1976_root_address, dout => ptr_deref_1976_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_267 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1976_base_resize_req_0;
      ptr_deref_1976_base_resize_ack_0 <= ack; 
      ptr_deref_1976_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep137_710, dout => ptr_deref_1976_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_268 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1980_addr_0_req_0;
      ptr_deref_1980_addr_0_ack_0 <= ack; 
      ptr_deref_1980_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1980_root_address, dout => ptr_deref_1980_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_269 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1980_base_resize_req_0;
      ptr_deref_1980_base_resize_ack_0 <= ack; 
      ptr_deref_1980_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep141_704, dout => ptr_deref_1980_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_270 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1984_addr_0_req_0;
      ptr_deref_1984_addr_0_ack_0 <= ack; 
      ptr_deref_1984_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1984_root_address, dout => ptr_deref_1984_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_271 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1984_base_resize_req_0;
      ptr_deref_1984_base_resize_ack_0 <= ack; 
      ptr_deref_1984_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep145_698, dout => ptr_deref_1984_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_272 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1988_addr_0_req_0;
      ptr_deref_1988_addr_0_ack_0 <= ack; 
      ptr_deref_1988_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1988_root_address, dout => ptr_deref_1988_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_273 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1988_base_resize_req_0;
      ptr_deref_1988_base_resize_ack_0 <= ack; 
      ptr_deref_1988_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep131_668, dout => ptr_deref_1988_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_274 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1992_addr_0_req_0;
      ptr_deref_1992_addr_0_ack_0 <= ack; 
      ptr_deref_1992_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1992_root_address, dout => ptr_deref_1992_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_275 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1992_base_resize_req_0;
      ptr_deref_1992_base_resize_ack_0 <= ack; 
      ptr_deref_1992_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep136_686, dout => ptr_deref_1992_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_276 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1996_addr_0_req_0;
      ptr_deref_1996_addr_0_ack_0 <= ack; 
      ptr_deref_1996_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_1996_root_address, dout => ptr_deref_1996_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_277 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_1996_base_resize_req_0;
      ptr_deref_1996_base_resize_ack_0 <= ack; 
      ptr_deref_1996_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep140_680, dout => ptr_deref_1996_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_278 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2000_addr_0_req_0;
      ptr_deref_2000_addr_0_ack_0 <= ack; 
      ptr_deref_2000_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_2000_root_address, dout => ptr_deref_2000_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_279 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2000_base_resize_req_0;
      ptr_deref_2000_base_resize_ack_0 <= ack; 
      ptr_deref_2000_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep144_674, dout => ptr_deref_2000_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_280 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2004_addr_0_req_0;
      ptr_deref_2004_addr_0_ack_0 <= ack; 
      ptr_deref_2004_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_2004_root_address, dout => ptr_deref_2004_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_281 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2004_base_resize_req_0;
      ptr_deref_2004_base_resize_ack_0 <= ack; 
      ptr_deref_2004_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep129_638, dout => ptr_deref_2004_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_282 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2008_addr_0_req_0;
      ptr_deref_2008_addr_0_ack_0 <= ack; 
      ptr_deref_2008_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_2008_root_address, dout => ptr_deref_2008_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_283 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2008_base_resize_req_0;
      ptr_deref_2008_base_resize_ack_0 <= ack; 
      ptr_deref_2008_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep135_662, dout => ptr_deref_2008_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_284 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2012_addr_0_req_0;
      ptr_deref_2012_addr_0_ack_0 <= ack; 
      ptr_deref_2012_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_2012_root_address, dout => ptr_deref_2012_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_285 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2012_base_resize_req_0;
      ptr_deref_2012_base_resize_ack_0 <= ack; 
      ptr_deref_2012_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep139_650, dout => ptr_deref_2012_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_286 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2016_addr_0_req_0;
      ptr_deref_2016_addr_0_ack_0 <= ack; 
      ptr_deref_2016_addr_0: RegisterBase --
        generic map(in_data_width => 9,out_data_width => 9) 
        port map( din => ptr_deref_2016_root_address, dout => ptr_deref_2016_word_address_0, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_287 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= ptr_deref_2016_base_resize_req_0;
      ptr_deref_2016_base_resize_ack_0 <= ack; 
      ptr_deref_2016_base_resize: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 9) 
        port map( din => scevgep143_644, dout => ptr_deref_2016_resized_base_address, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_288 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1893_inst_req_0;
      type_cast_1893_inst_ack_0 <= ack; 
      type_cast_1893_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_162_1870, dout => type_cast_1893_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_289 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1897_inst_req_0;
      type_cast_1897_inst_ack_0 <= ack; 
      type_cast_1897_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_154_1830, dout => type_cast_1897_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_290 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1901_inst_req_0;
      type_cast_1901_inst_ack_0 <= ack; 
      type_cast_1901_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_146_1790, dout => type_cast_1901_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_291 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1905_inst_req_0;
      type_cast_1905_inst_ack_0 <= ack; 
      type_cast_1905_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_138_1750, dout => type_cast_1905_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_292 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1909_inst_req_0;
      type_cast_1909_inst_ack_0 <= ack; 
      type_cast_1909_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_126_1694, dout => type_cast_1909_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_293 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1913_inst_req_0;
      type_cast_1913_inst_ack_0 <= ack; 
      type_cast_1913_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_118_1654, dout => type_cast_1913_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_294 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1917_inst_req_0;
      type_cast_1917_inst_ack_0 <= ack; 
      type_cast_1917_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_110_1614, dout => type_cast_1917_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_295 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1921_inst_req_0;
      type_cast_1921_inst_ack_0 <= ack; 
      type_cast_1921_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_102_1574, dout => type_cast_1921_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_296 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1925_inst_req_0;
      type_cast_1925_inst_ack_0 <= ack; 
      type_cast_1925_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_90_1518, dout => type_cast_1925_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_297 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1929_inst_req_0;
      type_cast_1929_inst_ack_0 <= ack; 
      type_cast_1929_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_82_1478, dout => type_cast_1929_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_298 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1933_inst_req_0;
      type_cast_1933_inst_ack_0 <= ack; 
      type_cast_1933_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_74_1438, dout => type_cast_1933_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_299 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1937_inst_req_0;
      type_cast_1937_inst_ack_0 <= ack; 
      type_cast_1937_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_66_1398, dout => type_cast_1937_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_300 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1941_inst_req_0;
      type_cast_1941_inst_ack_0 <= ack; 
      type_cast_1941_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_54_1342, dout => type_cast_1941_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_301 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1945_inst_req_0;
      type_cast_1945_inst_ack_0 <= ack; 
      type_cast_1945_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_42_1286, dout => type_cast_1945_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_302 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1949_inst_req_0;
      type_cast_1949_inst_ack_0 <= ack; 
      type_cast_1949_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_30_1230, dout => type_cast_1949_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_303 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1953_inst_req_0;
      type_cast_1953_inst_ack_0 <= ack; 
      type_cast_1953_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_18_1174, dout => type_cast_1953_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_304 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0 <= ack; 
      type_cast_561_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => indvarx_xnext61_2043, dout => type_cast_561_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_305 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_595_inst_req_0;
      type_cast_595_inst_ack_0 <= ack; 
      type_cast_595_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => indvarx_xnext57_2024, dout => type_cast_595_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_306 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_749_inst_req_0;
      type_cast_749_inst_ack_0 <= ack; 
      type_cast_749_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => indvarx_xnext_1876, dout => type_cast_749_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_307 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_756_inst_req_0;
      type_cast_756_inst_ack_0 <= ack; 
      type_cast_756_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_162_1870, dout => type_cast_756_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_308 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_763_inst_req_0;
      type_cast_763_inst_ack_0 <= ack; 
      type_cast_763_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_154_1830, dout => type_cast_763_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_309 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_770_inst_req_0;
      type_cast_770_inst_ack_0 <= ack; 
      type_cast_770_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_146_1790, dout => type_cast_770_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_310 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_777_inst_req_0;
      type_cast_777_inst_ack_0 <= ack; 
      type_cast_777_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_138_1750, dout => type_cast_777_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_311 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_784_inst_req_0;
      type_cast_784_inst_ack_0 <= ack; 
      type_cast_784_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_126_1694, dout => type_cast_784_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_312 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_791_inst_req_0;
      type_cast_791_inst_ack_0 <= ack; 
      type_cast_791_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_118_1654, dout => type_cast_791_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_313 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_798_inst_req_0;
      type_cast_798_inst_ack_0 <= ack; 
      type_cast_798_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_110_1614, dout => type_cast_798_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_314 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_805_inst_req_0;
      type_cast_805_inst_ack_0 <= ack; 
      type_cast_805_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_102_1574, dout => type_cast_805_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_315 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_812_inst_req_0;
      type_cast_812_inst_ack_0 <= ack; 
      type_cast_812_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_90_1518, dout => type_cast_812_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_316 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_819_inst_req_0;
      type_cast_819_inst_ack_0 <= ack; 
      type_cast_819_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_18_1174, dout => type_cast_819_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_317 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_826_inst_req_0;
      type_cast_826_inst_ack_0 <= ack; 
      type_cast_826_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_30_1230, dout => type_cast_826_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_318 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_833_inst_req_0;
      type_cast_833_inst_ack_0 <= ack; 
      type_cast_833_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_42_1286, dout => type_cast_833_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_319 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_840_inst_req_0;
      type_cast_840_inst_ack_0 <= ack; 
      type_cast_840_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_54_1342, dout => type_cast_840_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_320 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_847_inst_req_0;
      type_cast_847_inst_ack_0 <= ack; 
      type_cast_847_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_66_1398, dout => type_cast_847_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_321 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0 <= ack; 
      type_cast_854_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_74_1438, dout => type_cast_854_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    register_block_322 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_861_inst_req_0;
      type_cast_861_inst_ack_0 <= ack; 
      type_cast_861_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_82_1478, dout => type_cast_861_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    array_obj_ref_1010_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1010_index_1_rename_ack_0 <= array_obj_ref_1010_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1009_resized;
      simple_obj_ref_1009_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1010_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1010_root_address_inst_ack_0 <= array_obj_ref_1010_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1010_final_offset;
      array_obj_ref_1010_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1022_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1022_index_1_rename_ack_0 <= array_obj_ref_1022_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1021_resized;
      simple_obj_ref_1021_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1022_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1022_root_address_inst_ack_0 <= array_obj_ref_1022_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1022_final_offset;
      array_obj_ref_1022_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1028_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1028_index_1_rename_ack_0 <= array_obj_ref_1028_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1027_resized;
      simple_obj_ref_1027_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1028_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1028_root_address_inst_ack_0 <= array_obj_ref_1028_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1028_final_offset;
      array_obj_ref_1028_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1034_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1034_index_1_rename_ack_0 <= array_obj_ref_1034_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1033_resized;
      simple_obj_ref_1033_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1034_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1034_root_address_inst_ack_0 <= array_obj_ref_1034_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1034_final_offset;
      array_obj_ref_1034_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1040_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1040_index_1_rename_ack_0 <= array_obj_ref_1040_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1039_resized;
      simple_obj_ref_1039_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1040_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1040_root_address_inst_ack_0 <= array_obj_ref_1040_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1040_final_offset;
      array_obj_ref_1040_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1046_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1046_index_1_rename_ack_0 <= array_obj_ref_1046_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1045_resized;
      simple_obj_ref_1045_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1046_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1046_root_address_inst_ack_0 <= array_obj_ref_1046_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1046_final_offset;
      array_obj_ref_1046_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1052_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1052_index_1_rename_ack_0 <= array_obj_ref_1052_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1051_resized;
      simple_obj_ref_1051_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1052_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1052_root_address_inst_ack_0 <= array_obj_ref_1052_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1052_final_offset;
      array_obj_ref_1052_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1058_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1058_index_1_rename_ack_0 <= array_obj_ref_1058_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1057_resized;
      simple_obj_ref_1057_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1058_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1058_root_address_inst_ack_0 <= array_obj_ref_1058_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1058_final_offset;
      array_obj_ref_1058_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1064_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1064_index_1_rename_ack_0 <= array_obj_ref_1064_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1063_resized;
      simple_obj_ref_1063_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1064_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1064_root_address_inst_ack_0 <= array_obj_ref_1064_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1064_final_offset;
      array_obj_ref_1064_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1070_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1070_index_1_rename_ack_0 <= array_obj_ref_1070_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1069_resized;
      simple_obj_ref_1069_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1070_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1070_root_address_inst_ack_0 <= array_obj_ref_1070_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1070_final_offset;
      array_obj_ref_1070_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1076_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1076_index_1_rename_ack_0 <= array_obj_ref_1076_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1075_resized;
      simple_obj_ref_1075_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1076_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1076_root_address_inst_ack_0 <= array_obj_ref_1076_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1076_final_offset;
      array_obj_ref_1076_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1082_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1082_index_1_rename_ack_0 <= array_obj_ref_1082_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1081_resized;
      simple_obj_ref_1081_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1082_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1082_root_address_inst_ack_0 <= array_obj_ref_1082_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1082_final_offset;
      array_obj_ref_1082_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1088_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1088_index_1_rename_ack_0 <= array_obj_ref_1088_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1087_resized;
      simple_obj_ref_1087_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1088_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1088_root_address_inst_ack_0 <= array_obj_ref_1088_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1088_final_offset;
      array_obj_ref_1088_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1094_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1094_index_1_rename_ack_0 <= array_obj_ref_1094_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1093_resized;
      simple_obj_ref_1093_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1094_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1094_root_address_inst_ack_0 <= array_obj_ref_1094_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1094_final_offset;
      array_obj_ref_1094_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1100_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1100_index_1_rename_ack_0 <= array_obj_ref_1100_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_1099_resized;
      simple_obj_ref_1099_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_1100_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_1100_root_address_inst_ack_0 <= array_obj_ref_1100_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1100_final_offset;
      array_obj_ref_1100_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_606_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_606_index_1_rename_ack_0 <= array_obj_ref_606_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_605_resized;
      simple_obj_ref_605_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_606_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_606_root_address_inst_ack_0 <= array_obj_ref_606_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_606_final_offset;
      array_obj_ref_606_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_618_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_618_index_1_rename_ack_0 <= array_obj_ref_618_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_617_resized;
      simple_obj_ref_617_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_618_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_618_root_address_inst_ack_0 <= array_obj_ref_618_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_618_final_offset;
      array_obj_ref_618_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_630_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_630_index_1_rename_ack_0 <= array_obj_ref_630_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_629_resized;
      simple_obj_ref_629_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_630_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_630_root_address_inst_ack_0 <= array_obj_ref_630_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_630_final_offset;
      array_obj_ref_630_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_636_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_636_index_1_rename_ack_0 <= array_obj_ref_636_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_635_resized;
      simple_obj_ref_635_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_636_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_636_root_address_inst_ack_0 <= array_obj_ref_636_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_636_final_offset;
      array_obj_ref_636_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_642_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_642_index_1_rename_ack_0 <= array_obj_ref_642_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_641_resized;
      simple_obj_ref_641_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_642_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_642_root_address_inst_ack_0 <= array_obj_ref_642_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_642_final_offset;
      array_obj_ref_642_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_648_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_648_index_1_rename_ack_0 <= array_obj_ref_648_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_647_resized;
      simple_obj_ref_647_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_648_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_648_root_address_inst_ack_0 <= array_obj_ref_648_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_648_final_offset;
      array_obj_ref_648_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_660_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_660_index_1_rename_ack_0 <= array_obj_ref_660_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_659_resized;
      simple_obj_ref_659_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_660_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_660_root_address_inst_ack_0 <= array_obj_ref_660_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_660_final_offset;
      array_obj_ref_660_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_666_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_666_index_1_rename_ack_0 <= array_obj_ref_666_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_665_resized;
      simple_obj_ref_665_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_666_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_666_root_address_inst_ack_0 <= array_obj_ref_666_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_666_final_offset;
      array_obj_ref_666_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_672_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_672_index_1_rename_ack_0 <= array_obj_ref_672_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_671_resized;
      simple_obj_ref_671_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_672_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_672_root_address_inst_ack_0 <= array_obj_ref_672_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_672_final_offset;
      array_obj_ref_672_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_678_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_678_index_1_rename_ack_0 <= array_obj_ref_678_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_677_resized;
      simple_obj_ref_677_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_678_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_678_root_address_inst_ack_0 <= array_obj_ref_678_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_678_final_offset;
      array_obj_ref_678_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_684_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_684_index_1_rename_ack_0 <= array_obj_ref_684_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_683_resized;
      simple_obj_ref_683_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_684_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_684_root_address_inst_ack_0 <= array_obj_ref_684_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_684_final_offset;
      array_obj_ref_684_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_690_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_690_index_1_rename_ack_0 <= array_obj_ref_690_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_689_resized;
      simple_obj_ref_689_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_690_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_690_root_address_inst_ack_0 <= array_obj_ref_690_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_690_final_offset;
      array_obj_ref_690_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_696_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_696_index_1_rename_ack_0 <= array_obj_ref_696_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_695_resized;
      simple_obj_ref_695_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_696_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_696_root_address_inst_ack_0 <= array_obj_ref_696_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_696_final_offset;
      array_obj_ref_696_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_702_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_702_index_1_rename_ack_0 <= array_obj_ref_702_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_701_resized;
      simple_obj_ref_701_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_702_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_702_root_address_inst_ack_0 <= array_obj_ref_702_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_702_final_offset;
      array_obj_ref_702_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_708_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_708_index_1_rename_ack_0 <= array_obj_ref_708_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_707_resized;
      simple_obj_ref_707_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_708_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_708_root_address_inst_ack_0 <= array_obj_ref_708_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_708_final_offset;
      array_obj_ref_708_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_714_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_714_index_1_rename_ack_0 <= array_obj_ref_714_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_713_resized;
      simple_obj_ref_713_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_714_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_714_root_address_inst_ack_0 <= array_obj_ref_714_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_714_final_offset;
      array_obj_ref_714_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_872_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_872_index_1_rename_ack_0 <= array_obj_ref_872_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_871_resized;
      simple_obj_ref_871_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_872_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_872_root_address_inst_ack_0 <= array_obj_ref_872_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_872_final_offset;
      array_obj_ref_872_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_884_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_884_index_1_rename_ack_0 <= array_obj_ref_884_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_883_resized;
      simple_obj_ref_883_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_884_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_884_root_address_inst_ack_0 <= array_obj_ref_884_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_884_final_offset;
      array_obj_ref_884_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_896_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_896_index_1_rename_ack_0 <= array_obj_ref_896_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_895_resized;
      simple_obj_ref_895_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_896_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_896_root_address_inst_ack_0 <= array_obj_ref_896_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_896_final_offset;
      array_obj_ref_896_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_902_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_902_index_1_rename_ack_0 <= array_obj_ref_902_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_901_resized;
      simple_obj_ref_901_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_902_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_902_root_address_inst_ack_0 <= array_obj_ref_902_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_902_final_offset;
      array_obj_ref_902_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_908_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_908_index_1_rename_ack_0 <= array_obj_ref_908_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_907_resized;
      simple_obj_ref_907_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_908_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_908_root_address_inst_ack_0 <= array_obj_ref_908_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_908_final_offset;
      array_obj_ref_908_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_914_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_914_index_1_rename_ack_0 <= array_obj_ref_914_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_913_resized;
      simple_obj_ref_913_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_914_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_914_root_address_inst_ack_0 <= array_obj_ref_914_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_914_final_offset;
      array_obj_ref_914_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_926_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_926_index_1_rename_ack_0 <= array_obj_ref_926_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_925_resized;
      simple_obj_ref_925_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_926_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_926_root_address_inst_ack_0 <= array_obj_ref_926_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_926_final_offset;
      array_obj_ref_926_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_932_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_932_index_1_rename_ack_0 <= array_obj_ref_932_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_931_resized;
      simple_obj_ref_931_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_932_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_932_root_address_inst_ack_0 <= array_obj_ref_932_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_932_final_offset;
      array_obj_ref_932_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_938_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_938_index_1_rename_ack_0 <= array_obj_ref_938_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_937_resized;
      simple_obj_ref_937_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_938_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_938_root_address_inst_ack_0 <= array_obj_ref_938_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_938_final_offset;
      array_obj_ref_938_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_944_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_944_index_1_rename_ack_0 <= array_obj_ref_944_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_943_resized;
      simple_obj_ref_943_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_944_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_944_root_address_inst_ack_0 <= array_obj_ref_944_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_944_final_offset;
      array_obj_ref_944_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_950_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_950_index_1_rename_ack_0 <= array_obj_ref_950_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_949_resized;
      simple_obj_ref_949_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_950_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_950_root_address_inst_ack_0 <= array_obj_ref_950_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_950_final_offset;
      array_obj_ref_950_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_956_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_956_index_1_rename_ack_0 <= array_obj_ref_956_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_955_resized;
      simple_obj_ref_955_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_956_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_956_root_address_inst_ack_0 <= array_obj_ref_956_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_956_final_offset;
      array_obj_ref_956_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_962_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_962_index_1_rename_ack_0 <= array_obj_ref_962_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_961_resized;
      simple_obj_ref_961_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_962_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_962_root_address_inst_ack_0 <= array_obj_ref_962_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_962_final_offset;
      array_obj_ref_962_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_968_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_968_index_1_rename_ack_0 <= array_obj_ref_968_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_967_resized;
      simple_obj_ref_967_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_968_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_968_root_address_inst_ack_0 <= array_obj_ref_968_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_968_final_offset;
      array_obj_ref_968_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_974_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_974_index_1_rename_ack_0 <= array_obj_ref_974_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_973_resized;
      simple_obj_ref_973_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_974_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_974_root_address_inst_ack_0 <= array_obj_ref_974_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_974_final_offset;
      array_obj_ref_974_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_980_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_980_index_1_rename_ack_0 <= array_obj_ref_980_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_979_resized;
      simple_obj_ref_979_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_980_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_980_root_address_inst_ack_0 <= array_obj_ref_980_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_980_final_offset;
      array_obj_ref_980_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_998_index_1_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_998_index_1_rename_ack_0 <= array_obj_ref_998_index_1_rename_req_0;
      aggregated_sig <= simple_obj_ref_997_resized;
      simple_obj_ref_997_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_998_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_998_root_address_inst_ack_0 <= array_obj_ref_998_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_998_final_offset;
      array_obj_ref_998_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1105_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1105_gather_scatter_ack_0 <= ptr_deref_1105_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1105_data_0;
      iNsTr_3_1106 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1105_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1105_root_address_inst_ack_0 <= ptr_deref_1105_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1105_resized_base_address;
      ptr_deref_1105_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1109_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1109_gather_scatter_ack_0 <= ptr_deref_1109_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1109_data_0;
      iNsTr_4_1110 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1109_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1109_root_address_inst_ack_0 <= ptr_deref_1109_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1109_resized_base_address;
      ptr_deref_1109_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1113_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1113_gather_scatter_ack_0 <= ptr_deref_1113_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1113_data_0;
      iNsTr_5_1114 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1113_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1113_root_address_inst_ack_0 <= ptr_deref_1113_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1113_resized_base_address;
      ptr_deref_1113_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1117_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1117_gather_scatter_ack_0 <= ptr_deref_1117_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1117_data_0;
      iNsTr_6_1118 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1117_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1117_root_address_inst_ack_0 <= ptr_deref_1117_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1117_resized_base_address;
      ptr_deref_1117_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1121_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1121_gather_scatter_ack_0 <= ptr_deref_1121_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1121_data_0;
      iNsTr_7_1122 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1121_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1121_root_address_inst_ack_0 <= ptr_deref_1121_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1121_resized_base_address;
      ptr_deref_1121_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1125_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1125_gather_scatter_ack_0 <= ptr_deref_1125_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1125_data_0;
      iNsTr_8_1126 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1125_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1125_root_address_inst_ack_0 <= ptr_deref_1125_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1125_resized_base_address;
      ptr_deref_1125_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1129_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1129_gather_scatter_ack_0 <= ptr_deref_1129_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1129_data_0;
      iNsTr_9_1130 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1129_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1129_root_address_inst_ack_0 <= ptr_deref_1129_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1129_resized_base_address;
      ptr_deref_1129_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1133_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1133_gather_scatter_ack_0 <= ptr_deref_1133_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1133_data_0;
      iNsTr_10_1134 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1133_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1133_root_address_inst_ack_0 <= ptr_deref_1133_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1133_resized_base_address;
      ptr_deref_1133_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1177_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1177_gather_scatter_ack_0 <= ptr_deref_1177_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1177_data_0;
      iNsTr_19_1178 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1177_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1177_root_address_inst_ack_0 <= ptr_deref_1177_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1177_resized_base_address;
      ptr_deref_1177_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1181_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1181_gather_scatter_ack_0 <= ptr_deref_1181_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1181_data_0;
      iNsTr_20_1182 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1181_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1181_root_address_inst_ack_0 <= ptr_deref_1181_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1181_resized_base_address;
      ptr_deref_1181_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1185_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1185_gather_scatter_ack_0 <= ptr_deref_1185_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1185_data_0;
      iNsTr_21_1186 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1185_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1185_root_address_inst_ack_0 <= ptr_deref_1185_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1185_resized_base_address;
      ptr_deref_1185_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1189_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1189_gather_scatter_ack_0 <= ptr_deref_1189_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1189_data_0;
      iNsTr_22_1190 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1189_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1189_root_address_inst_ack_0 <= ptr_deref_1189_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1189_resized_base_address;
      ptr_deref_1189_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1233_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1233_gather_scatter_ack_0 <= ptr_deref_1233_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1233_data_0;
      iNsTr_31_1234 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1233_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1233_root_address_inst_ack_0 <= ptr_deref_1233_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1233_resized_base_address;
      ptr_deref_1233_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1237_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1237_gather_scatter_ack_0 <= ptr_deref_1237_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1237_data_0;
      iNsTr_32_1238 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1237_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1237_root_address_inst_ack_0 <= ptr_deref_1237_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1237_resized_base_address;
      ptr_deref_1237_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1241_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1241_gather_scatter_ack_0 <= ptr_deref_1241_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1241_data_0;
      iNsTr_33_1242 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1241_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1241_root_address_inst_ack_0 <= ptr_deref_1241_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1241_resized_base_address;
      ptr_deref_1241_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1245_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1245_gather_scatter_ack_0 <= ptr_deref_1245_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1245_data_0;
      iNsTr_34_1246 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1245_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1245_root_address_inst_ack_0 <= ptr_deref_1245_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1245_resized_base_address;
      ptr_deref_1245_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1289_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1289_gather_scatter_ack_0 <= ptr_deref_1289_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1289_data_0;
      iNsTr_43_1290 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1289_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1289_root_address_inst_ack_0 <= ptr_deref_1289_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1289_resized_base_address;
      ptr_deref_1289_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1293_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1293_gather_scatter_ack_0 <= ptr_deref_1293_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1293_data_0;
      iNsTr_44_1294 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1293_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1293_root_address_inst_ack_0 <= ptr_deref_1293_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1293_resized_base_address;
      ptr_deref_1293_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1297_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1297_gather_scatter_ack_0 <= ptr_deref_1297_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1297_data_0;
      iNsTr_45_1298 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1297_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1297_root_address_inst_ack_0 <= ptr_deref_1297_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1297_resized_base_address;
      ptr_deref_1297_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1301_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1301_gather_scatter_ack_0 <= ptr_deref_1301_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1301_data_0;
      iNsTr_46_1302 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1301_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1301_root_address_inst_ack_0 <= ptr_deref_1301_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1301_resized_base_address;
      ptr_deref_1301_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1345_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1345_gather_scatter_ack_0 <= ptr_deref_1345_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1345_data_0;
      iNsTr_55_1346 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1345_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1345_root_address_inst_ack_0 <= ptr_deref_1345_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1345_resized_base_address;
      ptr_deref_1345_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1349_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1349_gather_scatter_ack_0 <= ptr_deref_1349_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1349_data_0;
      iNsTr_56_1350 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1349_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1349_root_address_inst_ack_0 <= ptr_deref_1349_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1349_resized_base_address;
      ptr_deref_1349_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1353_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1353_gather_scatter_ack_0 <= ptr_deref_1353_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1353_data_0;
      iNsTr_57_1354 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1353_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1353_root_address_inst_ack_0 <= ptr_deref_1353_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1353_resized_base_address;
      ptr_deref_1353_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1357_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1357_gather_scatter_ack_0 <= ptr_deref_1357_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1357_data_0;
      iNsTr_58_1358 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1357_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1357_root_address_inst_ack_0 <= ptr_deref_1357_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1357_resized_base_address;
      ptr_deref_1357_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1521_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1521_gather_scatter_ack_0 <= ptr_deref_1521_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1521_data_0;
      iNsTr_91_1522 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1521_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1521_root_address_inst_ack_0 <= ptr_deref_1521_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1521_resized_base_address;
      ptr_deref_1521_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1525_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1525_gather_scatter_ack_0 <= ptr_deref_1525_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1525_data_0;
      iNsTr_92_1526 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1525_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1525_root_address_inst_ack_0 <= ptr_deref_1525_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1525_resized_base_address;
      ptr_deref_1525_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1529_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1529_gather_scatter_ack_0 <= ptr_deref_1529_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1529_data_0;
      iNsTr_93_1530 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1529_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1529_root_address_inst_ack_0 <= ptr_deref_1529_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1529_resized_base_address;
      ptr_deref_1529_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1533_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1533_gather_scatter_ack_0 <= ptr_deref_1533_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1533_data_0;
      iNsTr_94_1534 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1533_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1533_root_address_inst_ack_0 <= ptr_deref_1533_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1533_resized_base_address;
      ptr_deref_1533_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1697_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1697_gather_scatter_ack_0 <= ptr_deref_1697_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1697_data_0;
      iNsTr_127_1698 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1697_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1697_root_address_inst_ack_0 <= ptr_deref_1697_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1697_resized_base_address;
      ptr_deref_1697_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1701_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1701_gather_scatter_ack_0 <= ptr_deref_1701_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1701_data_0;
      iNsTr_128_1702 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1701_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1701_root_address_inst_ack_0 <= ptr_deref_1701_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1701_resized_base_address;
      ptr_deref_1701_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1705_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1705_gather_scatter_ack_0 <= ptr_deref_1705_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1705_data_0;
      iNsTr_129_1706 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1705_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1705_root_address_inst_ack_0 <= ptr_deref_1705_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1705_resized_base_address;
      ptr_deref_1705_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1709_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1709_gather_scatter_ack_0 <= ptr_deref_1709_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1709_data_0;
      iNsTr_130_1710 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1709_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1709_root_address_inst_ack_0 <= ptr_deref_1709_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1709_resized_base_address;
      ptr_deref_1709_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1956_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1956_gather_scatter_ack_0 <= ptr_deref_1956_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa_1950;
      ptr_deref_1956_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1956_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1956_root_address_inst_ack_0 <= ptr_deref_1956_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1956_resized_base_address;
      ptr_deref_1956_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1960_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1960_gather_scatter_ack_0 <= ptr_deref_1960_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa207_1946;
      ptr_deref_1960_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1960_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1960_root_address_inst_ack_0 <= ptr_deref_1960_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1960_resized_base_address;
      ptr_deref_1960_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1964_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1964_gather_scatter_ack_0 <= ptr_deref_1964_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa208_1942;
      ptr_deref_1964_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1964_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1964_root_address_inst_ack_0 <= ptr_deref_1964_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1964_resized_base_address;
      ptr_deref_1964_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1968_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1968_gather_scatter_ack_0 <= ptr_deref_1968_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa209_1938;
      ptr_deref_1968_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1968_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1968_root_address_inst_ack_0 <= ptr_deref_1968_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1968_resized_base_address;
      ptr_deref_1968_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1972_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1972_gather_scatter_ack_0 <= ptr_deref_1972_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa210_1934;
      ptr_deref_1972_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1972_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1972_root_address_inst_ack_0 <= ptr_deref_1972_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1972_resized_base_address;
      ptr_deref_1972_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1976_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1976_gather_scatter_ack_0 <= ptr_deref_1976_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa211_1930;
      ptr_deref_1976_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1976_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1976_root_address_inst_ack_0 <= ptr_deref_1976_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1976_resized_base_address;
      ptr_deref_1976_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1980_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1980_gather_scatter_ack_0 <= ptr_deref_1980_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa212_1926;
      ptr_deref_1980_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1980_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1980_root_address_inst_ack_0 <= ptr_deref_1980_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1980_resized_base_address;
      ptr_deref_1980_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1984_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1984_gather_scatter_ack_0 <= ptr_deref_1984_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa213_1922;
      ptr_deref_1984_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1984_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1984_root_address_inst_ack_0 <= ptr_deref_1984_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1984_resized_base_address;
      ptr_deref_1984_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1988_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1988_gather_scatter_ack_0 <= ptr_deref_1988_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa214_1918;
      ptr_deref_1988_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1988_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1988_root_address_inst_ack_0 <= ptr_deref_1988_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1988_resized_base_address;
      ptr_deref_1988_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1992_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1992_gather_scatter_ack_0 <= ptr_deref_1992_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa215_1914;
      ptr_deref_1992_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1992_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1992_root_address_inst_ack_0 <= ptr_deref_1992_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1992_resized_base_address;
      ptr_deref_1992_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1996_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1996_gather_scatter_ack_0 <= ptr_deref_1996_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa216_1910;
      ptr_deref_1996_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1996_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_1996_root_address_inst_ack_0 <= ptr_deref_1996_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1996_resized_base_address;
      ptr_deref_1996_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2000_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2000_gather_scatter_ack_0 <= ptr_deref_2000_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa217_1906;
      ptr_deref_2000_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2000_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2000_root_address_inst_ack_0 <= ptr_deref_2000_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2000_resized_base_address;
      ptr_deref_2000_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2004_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2004_gather_scatter_ack_0 <= ptr_deref_2004_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa218_1902;
      ptr_deref_2004_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2004_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2004_root_address_inst_ack_0 <= ptr_deref_2004_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2004_resized_base_address;
      ptr_deref_2004_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2008_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2008_gather_scatter_ack_0 <= ptr_deref_2008_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa219_1898;
      ptr_deref_2008_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2008_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2008_root_address_inst_ack_0 <= ptr_deref_2008_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2008_resized_base_address;
      ptr_deref_2008_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2012_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2012_gather_scatter_ack_0 <= ptr_deref_2012_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa220_1894;
      ptr_deref_2012_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2012_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2012_root_address_inst_ack_0 <= ptr_deref_2012_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2012_resized_base_address;
      ptr_deref_2012_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2016_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2016_gather_scatter_ack_0 <= ptr_deref_2016_gather_scatter_req_0;
      aggregated_sig <= xx_xlcssa221_1890;
      ptr_deref_2016_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2016_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2016_root_address_inst_ack_0 <= ptr_deref_2016_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2016_resized_base_address;
      ptr_deref_2016_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    if_stmt_1883_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond222_1882;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1883_branch_req_0,
          ack0 => if_stmt_1883_branch_ack_0,
          ack1 => if_stmt_1883_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2031_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_2030;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2031_branch_req_0,
          ack0 => if_stmt_2031_branch_ack_0,
          ack1 => if_stmt_2031_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2050_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond310_2049;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2050_branch_req_0,
          ack0 => if_stmt_2050_branch_ack_0,
          ack1 => if_stmt_2050_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_950_index_0_scale array_obj_ref_944_index_0_scale array_obj_ref_980_index_0_scale array_obj_ref_938_index_0_scale array_obj_ref_926_index_0_scale array_obj_ref_974_index_0_scale array_obj_ref_956_index_0_scale array_obj_ref_1028_index_0_scale array_obj_ref_914_index_0_scale array_obj_ref_1022_index_0_scale array_obj_ref_932_index_0_scale array_obj_ref_1034_index_0_scale array_obj_ref_1040_index_0_scale array_obj_ref_998_index_0_scale array_obj_ref_908_index_0_scale array_obj_ref_1076_index_0_scale array_obj_ref_962_index_0_scale array_obj_ref_1064_index_0_scale array_obj_ref_1070_index_0_scale array_obj_ref_1052_index_0_scale array_obj_ref_1046_index_0_scale array_obj_ref_968_index_0_scale array_obj_ref_1058_index_0_scale array_obj_ref_1010_index_0_scale array_obj_ref_902_index_0_scale array_obj_ref_896_index_0_scale array_obj_ref_1082_index_0_scale array_obj_ref_1094_index_0_scale array_obj_ref_872_index_0_scale array_obj_ref_884_index_0_scale array_obj_ref_1088_index_0_scale array_obj_ref_606_index_0_scale array_obj_ref_618_index_0_scale array_obj_ref_630_index_0_scale array_obj_ref_636_index_0_scale array_obj_ref_642_index_0_scale array_obj_ref_648_index_0_scale array_obj_ref_660_index_0_scale array_obj_ref_666_index_0_scale array_obj_ref_672_index_0_scale array_obj_ref_678_index_0_scale array_obj_ref_684_index_0_scale array_obj_ref_690_index_0_scale array_obj_ref_696_index_0_scale array_obj_ref_702_index_0_scale array_obj_ref_708_index_0_scale array_obj_ref_714_index_0_scale array_obj_ref_1100_index_0_scale 
    ApIntMul_group_0: Block -- 
      signal data_in: std_logic_vector(431 downto 0);
      signal data_out: std_logic_vector(431 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 47 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 47 downto 0);
      signal guard_vector : std_logic_vector( 47 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_948_resized & simple_obj_ref_942_resized & simple_obj_ref_978_resized & simple_obj_ref_936_resized & simple_obj_ref_924_resized & simple_obj_ref_972_resized & simple_obj_ref_954_resized & simple_obj_ref_1026_resized & simple_obj_ref_912_resized & simple_obj_ref_1020_resized & simple_obj_ref_930_resized & simple_obj_ref_1032_resized & simple_obj_ref_1038_resized & simple_obj_ref_996_resized & simple_obj_ref_906_resized & simple_obj_ref_1074_resized & simple_obj_ref_960_resized & simple_obj_ref_1062_resized & simple_obj_ref_1068_resized & simple_obj_ref_1050_resized & simple_obj_ref_1044_resized & simple_obj_ref_966_resized & simple_obj_ref_1056_resized & simple_obj_ref_1008_resized & simple_obj_ref_900_resized & simple_obj_ref_894_resized & simple_obj_ref_1080_resized & simple_obj_ref_1092_resized & simple_obj_ref_870_resized & simple_obj_ref_882_resized & simple_obj_ref_1086_resized & simple_obj_ref_604_resized & simple_obj_ref_616_resized & simple_obj_ref_628_resized & simple_obj_ref_634_resized & simple_obj_ref_640_resized & simple_obj_ref_646_resized & simple_obj_ref_658_resized & simple_obj_ref_664_resized & simple_obj_ref_670_resized & simple_obj_ref_676_resized & simple_obj_ref_682_resized & simple_obj_ref_688_resized & simple_obj_ref_694_resized & simple_obj_ref_700_resized & simple_obj_ref_706_resized & simple_obj_ref_712_resized & simple_obj_ref_1098_resized;
      simple_obj_ref_948_scaled <= data_out(431 downto 423);
      simple_obj_ref_942_scaled <= data_out(422 downto 414);
      simple_obj_ref_978_scaled <= data_out(413 downto 405);
      simple_obj_ref_936_scaled <= data_out(404 downto 396);
      simple_obj_ref_924_scaled <= data_out(395 downto 387);
      simple_obj_ref_972_scaled <= data_out(386 downto 378);
      simple_obj_ref_954_scaled <= data_out(377 downto 369);
      simple_obj_ref_1026_scaled <= data_out(368 downto 360);
      simple_obj_ref_912_scaled <= data_out(359 downto 351);
      simple_obj_ref_1020_scaled <= data_out(350 downto 342);
      simple_obj_ref_930_scaled <= data_out(341 downto 333);
      simple_obj_ref_1032_scaled <= data_out(332 downto 324);
      simple_obj_ref_1038_scaled <= data_out(323 downto 315);
      simple_obj_ref_996_scaled <= data_out(314 downto 306);
      simple_obj_ref_906_scaled <= data_out(305 downto 297);
      simple_obj_ref_1074_scaled <= data_out(296 downto 288);
      simple_obj_ref_960_scaled <= data_out(287 downto 279);
      simple_obj_ref_1062_scaled <= data_out(278 downto 270);
      simple_obj_ref_1068_scaled <= data_out(269 downto 261);
      simple_obj_ref_1050_scaled <= data_out(260 downto 252);
      simple_obj_ref_1044_scaled <= data_out(251 downto 243);
      simple_obj_ref_966_scaled <= data_out(242 downto 234);
      simple_obj_ref_1056_scaled <= data_out(233 downto 225);
      simple_obj_ref_1008_scaled <= data_out(224 downto 216);
      simple_obj_ref_900_scaled <= data_out(215 downto 207);
      simple_obj_ref_894_scaled <= data_out(206 downto 198);
      simple_obj_ref_1080_scaled <= data_out(197 downto 189);
      simple_obj_ref_1092_scaled <= data_out(188 downto 180);
      simple_obj_ref_870_scaled <= data_out(179 downto 171);
      simple_obj_ref_882_scaled <= data_out(170 downto 162);
      simple_obj_ref_1086_scaled <= data_out(161 downto 153);
      simple_obj_ref_604_scaled <= data_out(152 downto 144);
      simple_obj_ref_616_scaled <= data_out(143 downto 135);
      simple_obj_ref_628_scaled <= data_out(134 downto 126);
      simple_obj_ref_634_scaled <= data_out(125 downto 117);
      simple_obj_ref_640_scaled <= data_out(116 downto 108);
      simple_obj_ref_646_scaled <= data_out(107 downto 99);
      simple_obj_ref_658_scaled <= data_out(98 downto 90);
      simple_obj_ref_664_scaled <= data_out(89 downto 81);
      simple_obj_ref_670_scaled <= data_out(80 downto 72);
      simple_obj_ref_676_scaled <= data_out(71 downto 63);
      simple_obj_ref_682_scaled <= data_out(62 downto 54);
      simple_obj_ref_688_scaled <= data_out(53 downto 45);
      simple_obj_ref_694_scaled <= data_out(44 downto 36);
      simple_obj_ref_700_scaled <= data_out(35 downto 27);
      simple_obj_ref_706_scaled <= data_out(26 downto 18);
      simple_obj_ref_712_scaled <= data_out(17 downto 9);
      simple_obj_ref_1098_scaled <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      guard_vector(40)  <=  '1';
      guard_vector(41)  <=  '1';
      guard_vector(42)  <=  '1';
      guard_vector(43)  <=  '1';
      guard_vector(44)  <=  '1';
      guard_vector(45)  <=  '1';
      guard_vector(46)  <=  '1';
      guard_vector(47)  <=  '1';
      reqL_unguarded(47) <= array_obj_ref_950_index_0_scale_req_0;
      reqL_unguarded(46) <= array_obj_ref_944_index_0_scale_req_0;
      reqL_unguarded(45) <= array_obj_ref_980_index_0_scale_req_0;
      reqL_unguarded(44) <= array_obj_ref_938_index_0_scale_req_0;
      reqL_unguarded(43) <= array_obj_ref_926_index_0_scale_req_0;
      reqL_unguarded(42) <= array_obj_ref_974_index_0_scale_req_0;
      reqL_unguarded(41) <= array_obj_ref_956_index_0_scale_req_0;
      reqL_unguarded(40) <= array_obj_ref_1028_index_0_scale_req_0;
      reqL_unguarded(39) <= array_obj_ref_914_index_0_scale_req_0;
      reqL_unguarded(38) <= array_obj_ref_1022_index_0_scale_req_0;
      reqL_unguarded(37) <= array_obj_ref_932_index_0_scale_req_0;
      reqL_unguarded(36) <= array_obj_ref_1034_index_0_scale_req_0;
      reqL_unguarded(35) <= array_obj_ref_1040_index_0_scale_req_0;
      reqL_unguarded(34) <= array_obj_ref_998_index_0_scale_req_0;
      reqL_unguarded(33) <= array_obj_ref_908_index_0_scale_req_0;
      reqL_unguarded(32) <= array_obj_ref_1076_index_0_scale_req_0;
      reqL_unguarded(31) <= array_obj_ref_962_index_0_scale_req_0;
      reqL_unguarded(30) <= array_obj_ref_1064_index_0_scale_req_0;
      reqL_unguarded(29) <= array_obj_ref_1070_index_0_scale_req_0;
      reqL_unguarded(28) <= array_obj_ref_1052_index_0_scale_req_0;
      reqL_unguarded(27) <= array_obj_ref_1046_index_0_scale_req_0;
      reqL_unguarded(26) <= array_obj_ref_968_index_0_scale_req_0;
      reqL_unguarded(25) <= array_obj_ref_1058_index_0_scale_req_0;
      reqL_unguarded(24) <= array_obj_ref_1010_index_0_scale_req_0;
      reqL_unguarded(23) <= array_obj_ref_902_index_0_scale_req_0;
      reqL_unguarded(22) <= array_obj_ref_896_index_0_scale_req_0;
      reqL_unguarded(21) <= array_obj_ref_1082_index_0_scale_req_0;
      reqL_unguarded(20) <= array_obj_ref_1094_index_0_scale_req_0;
      reqL_unguarded(19) <= array_obj_ref_872_index_0_scale_req_0;
      reqL_unguarded(18) <= array_obj_ref_884_index_0_scale_req_0;
      reqL_unguarded(17) <= array_obj_ref_1088_index_0_scale_req_0;
      reqL_unguarded(16) <= array_obj_ref_606_index_0_scale_req_0;
      reqL_unguarded(15) <= array_obj_ref_618_index_0_scale_req_0;
      reqL_unguarded(14) <= array_obj_ref_630_index_0_scale_req_0;
      reqL_unguarded(13) <= array_obj_ref_636_index_0_scale_req_0;
      reqL_unguarded(12) <= array_obj_ref_642_index_0_scale_req_0;
      reqL_unguarded(11) <= array_obj_ref_648_index_0_scale_req_0;
      reqL_unguarded(10) <= array_obj_ref_660_index_0_scale_req_0;
      reqL_unguarded(9) <= array_obj_ref_666_index_0_scale_req_0;
      reqL_unguarded(8) <= array_obj_ref_672_index_0_scale_req_0;
      reqL_unguarded(7) <= array_obj_ref_678_index_0_scale_req_0;
      reqL_unguarded(6) <= array_obj_ref_684_index_0_scale_req_0;
      reqL_unguarded(5) <= array_obj_ref_690_index_0_scale_req_0;
      reqL_unguarded(4) <= array_obj_ref_696_index_0_scale_req_0;
      reqL_unguarded(3) <= array_obj_ref_702_index_0_scale_req_0;
      reqL_unguarded(2) <= array_obj_ref_708_index_0_scale_req_0;
      reqL_unguarded(1) <= array_obj_ref_714_index_0_scale_req_0;
      reqL_unguarded(0) <= array_obj_ref_1100_index_0_scale_req_0;
      array_obj_ref_950_index_0_scale_ack_0 <= ackL_unguarded(47);
      array_obj_ref_944_index_0_scale_ack_0 <= ackL_unguarded(46);
      array_obj_ref_980_index_0_scale_ack_0 <= ackL_unguarded(45);
      array_obj_ref_938_index_0_scale_ack_0 <= ackL_unguarded(44);
      array_obj_ref_926_index_0_scale_ack_0 <= ackL_unguarded(43);
      array_obj_ref_974_index_0_scale_ack_0 <= ackL_unguarded(42);
      array_obj_ref_956_index_0_scale_ack_0 <= ackL_unguarded(41);
      array_obj_ref_1028_index_0_scale_ack_0 <= ackL_unguarded(40);
      array_obj_ref_914_index_0_scale_ack_0 <= ackL_unguarded(39);
      array_obj_ref_1022_index_0_scale_ack_0 <= ackL_unguarded(38);
      array_obj_ref_932_index_0_scale_ack_0 <= ackL_unguarded(37);
      array_obj_ref_1034_index_0_scale_ack_0 <= ackL_unguarded(36);
      array_obj_ref_1040_index_0_scale_ack_0 <= ackL_unguarded(35);
      array_obj_ref_998_index_0_scale_ack_0 <= ackL_unguarded(34);
      array_obj_ref_908_index_0_scale_ack_0 <= ackL_unguarded(33);
      array_obj_ref_1076_index_0_scale_ack_0 <= ackL_unguarded(32);
      array_obj_ref_962_index_0_scale_ack_0 <= ackL_unguarded(31);
      array_obj_ref_1064_index_0_scale_ack_0 <= ackL_unguarded(30);
      array_obj_ref_1070_index_0_scale_ack_0 <= ackL_unguarded(29);
      array_obj_ref_1052_index_0_scale_ack_0 <= ackL_unguarded(28);
      array_obj_ref_1046_index_0_scale_ack_0 <= ackL_unguarded(27);
      array_obj_ref_968_index_0_scale_ack_0 <= ackL_unguarded(26);
      array_obj_ref_1058_index_0_scale_ack_0 <= ackL_unguarded(25);
      array_obj_ref_1010_index_0_scale_ack_0 <= ackL_unguarded(24);
      array_obj_ref_902_index_0_scale_ack_0 <= ackL_unguarded(23);
      array_obj_ref_896_index_0_scale_ack_0 <= ackL_unguarded(22);
      array_obj_ref_1082_index_0_scale_ack_0 <= ackL_unguarded(21);
      array_obj_ref_1094_index_0_scale_ack_0 <= ackL_unguarded(20);
      array_obj_ref_872_index_0_scale_ack_0 <= ackL_unguarded(19);
      array_obj_ref_884_index_0_scale_ack_0 <= ackL_unguarded(18);
      array_obj_ref_1088_index_0_scale_ack_0 <= ackL_unguarded(17);
      array_obj_ref_606_index_0_scale_ack_0 <= ackL_unguarded(16);
      array_obj_ref_618_index_0_scale_ack_0 <= ackL_unguarded(15);
      array_obj_ref_630_index_0_scale_ack_0 <= ackL_unguarded(14);
      array_obj_ref_636_index_0_scale_ack_0 <= ackL_unguarded(13);
      array_obj_ref_642_index_0_scale_ack_0 <= ackL_unguarded(12);
      array_obj_ref_648_index_0_scale_ack_0 <= ackL_unguarded(11);
      array_obj_ref_660_index_0_scale_ack_0 <= ackL_unguarded(10);
      array_obj_ref_666_index_0_scale_ack_0 <= ackL_unguarded(9);
      array_obj_ref_672_index_0_scale_ack_0 <= ackL_unguarded(8);
      array_obj_ref_678_index_0_scale_ack_0 <= ackL_unguarded(7);
      array_obj_ref_684_index_0_scale_ack_0 <= ackL_unguarded(6);
      array_obj_ref_690_index_0_scale_ack_0 <= ackL_unguarded(5);
      array_obj_ref_696_index_0_scale_ack_0 <= ackL_unguarded(4);
      array_obj_ref_702_index_0_scale_ack_0 <= ackL_unguarded(3);
      array_obj_ref_708_index_0_scale_ack_0 <= ackL_unguarded(2);
      array_obj_ref_714_index_0_scale_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1100_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(47) <= array_obj_ref_950_index_0_scale_req_1;
      reqR_unguarded(46) <= array_obj_ref_944_index_0_scale_req_1;
      reqR_unguarded(45) <= array_obj_ref_980_index_0_scale_req_1;
      reqR_unguarded(44) <= array_obj_ref_938_index_0_scale_req_1;
      reqR_unguarded(43) <= array_obj_ref_926_index_0_scale_req_1;
      reqR_unguarded(42) <= array_obj_ref_974_index_0_scale_req_1;
      reqR_unguarded(41) <= array_obj_ref_956_index_0_scale_req_1;
      reqR_unguarded(40) <= array_obj_ref_1028_index_0_scale_req_1;
      reqR_unguarded(39) <= array_obj_ref_914_index_0_scale_req_1;
      reqR_unguarded(38) <= array_obj_ref_1022_index_0_scale_req_1;
      reqR_unguarded(37) <= array_obj_ref_932_index_0_scale_req_1;
      reqR_unguarded(36) <= array_obj_ref_1034_index_0_scale_req_1;
      reqR_unguarded(35) <= array_obj_ref_1040_index_0_scale_req_1;
      reqR_unguarded(34) <= array_obj_ref_998_index_0_scale_req_1;
      reqR_unguarded(33) <= array_obj_ref_908_index_0_scale_req_1;
      reqR_unguarded(32) <= array_obj_ref_1076_index_0_scale_req_1;
      reqR_unguarded(31) <= array_obj_ref_962_index_0_scale_req_1;
      reqR_unguarded(30) <= array_obj_ref_1064_index_0_scale_req_1;
      reqR_unguarded(29) <= array_obj_ref_1070_index_0_scale_req_1;
      reqR_unguarded(28) <= array_obj_ref_1052_index_0_scale_req_1;
      reqR_unguarded(27) <= array_obj_ref_1046_index_0_scale_req_1;
      reqR_unguarded(26) <= array_obj_ref_968_index_0_scale_req_1;
      reqR_unguarded(25) <= array_obj_ref_1058_index_0_scale_req_1;
      reqR_unguarded(24) <= array_obj_ref_1010_index_0_scale_req_1;
      reqR_unguarded(23) <= array_obj_ref_902_index_0_scale_req_1;
      reqR_unguarded(22) <= array_obj_ref_896_index_0_scale_req_1;
      reqR_unguarded(21) <= array_obj_ref_1082_index_0_scale_req_1;
      reqR_unguarded(20) <= array_obj_ref_1094_index_0_scale_req_1;
      reqR_unguarded(19) <= array_obj_ref_872_index_0_scale_req_1;
      reqR_unguarded(18) <= array_obj_ref_884_index_0_scale_req_1;
      reqR_unguarded(17) <= array_obj_ref_1088_index_0_scale_req_1;
      reqR_unguarded(16) <= array_obj_ref_606_index_0_scale_req_1;
      reqR_unguarded(15) <= array_obj_ref_618_index_0_scale_req_1;
      reqR_unguarded(14) <= array_obj_ref_630_index_0_scale_req_1;
      reqR_unguarded(13) <= array_obj_ref_636_index_0_scale_req_1;
      reqR_unguarded(12) <= array_obj_ref_642_index_0_scale_req_1;
      reqR_unguarded(11) <= array_obj_ref_648_index_0_scale_req_1;
      reqR_unguarded(10) <= array_obj_ref_660_index_0_scale_req_1;
      reqR_unguarded(9) <= array_obj_ref_666_index_0_scale_req_1;
      reqR_unguarded(8) <= array_obj_ref_672_index_0_scale_req_1;
      reqR_unguarded(7) <= array_obj_ref_678_index_0_scale_req_1;
      reqR_unguarded(6) <= array_obj_ref_684_index_0_scale_req_1;
      reqR_unguarded(5) <= array_obj_ref_690_index_0_scale_req_1;
      reqR_unguarded(4) <= array_obj_ref_696_index_0_scale_req_1;
      reqR_unguarded(3) <= array_obj_ref_702_index_0_scale_req_1;
      reqR_unguarded(2) <= array_obj_ref_708_index_0_scale_req_1;
      reqR_unguarded(1) <= array_obj_ref_714_index_0_scale_req_1;
      reqR_unguarded(0) <= array_obj_ref_1100_index_0_scale_req_1;
      array_obj_ref_950_index_0_scale_ack_1 <= ackR_unguarded(47);
      array_obj_ref_944_index_0_scale_ack_1 <= ackR_unguarded(46);
      array_obj_ref_980_index_0_scale_ack_1 <= ackR_unguarded(45);
      array_obj_ref_938_index_0_scale_ack_1 <= ackR_unguarded(44);
      array_obj_ref_926_index_0_scale_ack_1 <= ackR_unguarded(43);
      array_obj_ref_974_index_0_scale_ack_1 <= ackR_unguarded(42);
      array_obj_ref_956_index_0_scale_ack_1 <= ackR_unguarded(41);
      array_obj_ref_1028_index_0_scale_ack_1 <= ackR_unguarded(40);
      array_obj_ref_914_index_0_scale_ack_1 <= ackR_unguarded(39);
      array_obj_ref_1022_index_0_scale_ack_1 <= ackR_unguarded(38);
      array_obj_ref_932_index_0_scale_ack_1 <= ackR_unguarded(37);
      array_obj_ref_1034_index_0_scale_ack_1 <= ackR_unguarded(36);
      array_obj_ref_1040_index_0_scale_ack_1 <= ackR_unguarded(35);
      array_obj_ref_998_index_0_scale_ack_1 <= ackR_unguarded(34);
      array_obj_ref_908_index_0_scale_ack_1 <= ackR_unguarded(33);
      array_obj_ref_1076_index_0_scale_ack_1 <= ackR_unguarded(32);
      array_obj_ref_962_index_0_scale_ack_1 <= ackR_unguarded(31);
      array_obj_ref_1064_index_0_scale_ack_1 <= ackR_unguarded(30);
      array_obj_ref_1070_index_0_scale_ack_1 <= ackR_unguarded(29);
      array_obj_ref_1052_index_0_scale_ack_1 <= ackR_unguarded(28);
      array_obj_ref_1046_index_0_scale_ack_1 <= ackR_unguarded(27);
      array_obj_ref_968_index_0_scale_ack_1 <= ackR_unguarded(26);
      array_obj_ref_1058_index_0_scale_ack_1 <= ackR_unguarded(25);
      array_obj_ref_1010_index_0_scale_ack_1 <= ackR_unguarded(24);
      array_obj_ref_902_index_0_scale_ack_1 <= ackR_unguarded(23);
      array_obj_ref_896_index_0_scale_ack_1 <= ackR_unguarded(22);
      array_obj_ref_1082_index_0_scale_ack_1 <= ackR_unguarded(21);
      array_obj_ref_1094_index_0_scale_ack_1 <= ackR_unguarded(20);
      array_obj_ref_872_index_0_scale_ack_1 <= ackR_unguarded(19);
      array_obj_ref_884_index_0_scale_ack_1 <= ackR_unguarded(18);
      array_obj_ref_1088_index_0_scale_ack_1 <= ackR_unguarded(17);
      array_obj_ref_606_index_0_scale_ack_1 <= ackR_unguarded(16);
      array_obj_ref_618_index_0_scale_ack_1 <= ackR_unguarded(15);
      array_obj_ref_630_index_0_scale_ack_1 <= ackR_unguarded(14);
      array_obj_ref_636_index_0_scale_ack_1 <= ackR_unguarded(13);
      array_obj_ref_642_index_0_scale_ack_1 <= ackR_unguarded(12);
      array_obj_ref_648_index_0_scale_ack_1 <= ackR_unguarded(11);
      array_obj_ref_660_index_0_scale_ack_1 <= ackR_unguarded(10);
      array_obj_ref_666_index_0_scale_ack_1 <= ackR_unguarded(9);
      array_obj_ref_672_index_0_scale_ack_1 <= ackR_unguarded(8);
      array_obj_ref_678_index_0_scale_ack_1 <= ackR_unguarded(7);
      array_obj_ref_684_index_0_scale_ack_1 <= ackR_unguarded(6);
      array_obj_ref_690_index_0_scale_ack_1 <= ackR_unguarded(5);
      array_obj_ref_696_index_0_scale_ack_1 <= ackR_unguarded(4);
      array_obj_ref_702_index_0_scale_ack_1 <= ackR_unguarded(3);
      array_obj_ref_708_index_0_scale_ack_1 <= ackR_unguarded(2);
      array_obj_ref_714_index_0_scale_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1100_index_0_scale_ack_1 <= ackR_unguarded(0);
      gI0: GuardInterface generic map(nreqs => 48) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 48) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000010000",
          constant_width => 9,
          use_constant  => true,
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 48--
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1010_index_sum_1 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1009_scaled & simple_obj_ref_1008_scaled;
      array_obj_ref_1010_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1010_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1010_index_sum_1_req_1;
      array_obj_ref_1010_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1010_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1022_index_sum_1 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1021_scaled & simple_obj_ref_1020_scaled;
      array_obj_ref_1022_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1022_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1022_index_sum_1_req_1;
      array_obj_ref_1022_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1022_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1028_index_sum_1 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1027_scaled & simple_obj_ref_1026_scaled;
      array_obj_ref_1028_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1028_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1028_index_sum_1_req_1;
      array_obj_ref_1028_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1028_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1034_index_sum_1 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1033_scaled & simple_obj_ref_1032_scaled;
      array_obj_ref_1034_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1034_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1034_index_sum_1_req_1;
      array_obj_ref_1034_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1034_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1040_index_sum_1 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1039_scaled & simple_obj_ref_1038_scaled;
      array_obj_ref_1040_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1040_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1040_index_sum_1_req_1;
      array_obj_ref_1040_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1040_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1046_index_sum_1 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1045_scaled & simple_obj_ref_1044_scaled;
      array_obj_ref_1046_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1046_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1046_index_sum_1_req_1;
      array_obj_ref_1046_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1046_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_1052_index_sum_1 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1051_scaled & simple_obj_ref_1050_scaled;
      array_obj_ref_1052_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1052_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1052_index_sum_1_req_1;
      array_obj_ref_1052_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1052_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_1058_index_sum_1 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1057_scaled & simple_obj_ref_1056_scaled;
      array_obj_ref_1058_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1058_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1058_index_sum_1_req_1;
      array_obj_ref_1058_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1058_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_1064_index_sum_1 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1063_scaled & simple_obj_ref_1062_scaled;
      array_obj_ref_1064_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1064_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1064_index_sum_1_req_1;
      array_obj_ref_1064_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1064_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_1070_index_sum_1 
    ApIntAdd_group_10: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1069_scaled & simple_obj_ref_1068_scaled;
      array_obj_ref_1070_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1070_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1070_index_sum_1_req_1;
      array_obj_ref_1070_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1070_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_1076_index_sum_1 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1075_scaled & simple_obj_ref_1074_scaled;
      array_obj_ref_1076_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1076_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1076_index_sum_1_req_1;
      array_obj_ref_1076_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1076_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_1082_index_sum_1 
    ApIntAdd_group_12: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1081_scaled & simple_obj_ref_1080_scaled;
      array_obj_ref_1082_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1082_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1082_index_sum_1_req_1;
      array_obj_ref_1082_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1082_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_1088_index_sum_1 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1087_scaled & simple_obj_ref_1086_scaled;
      array_obj_ref_1088_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1088_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1088_index_sum_1_req_1;
      array_obj_ref_1088_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1088_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_1094_index_sum_1 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1093_scaled & simple_obj_ref_1092_scaled;
      array_obj_ref_1094_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1094_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1094_index_sum_1_req_1;
      array_obj_ref_1094_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1094_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : array_obj_ref_1100_index_sum_1 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1099_scaled & simple_obj_ref_1098_scaled;
      array_obj_ref_1100_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_1100_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_1100_index_sum_1_req_1;
      array_obj_ref_1100_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_1100_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : array_obj_ref_606_index_sum_1 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_605_scaled & simple_obj_ref_604_scaled;
      array_obj_ref_606_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_606_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_606_index_sum_1_req_1;
      array_obj_ref_606_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_606_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : array_obj_ref_618_index_sum_1 
    ApIntAdd_group_17: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_617_scaled & simple_obj_ref_616_scaled;
      array_obj_ref_618_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_618_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_618_index_sum_1_req_1;
      array_obj_ref_618_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_618_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : array_obj_ref_630_index_sum_1 
    ApIntAdd_group_18: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_629_scaled & simple_obj_ref_628_scaled;
      array_obj_ref_630_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_630_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_630_index_sum_1_req_1;
      array_obj_ref_630_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_630_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : array_obj_ref_636_index_sum_1 
    ApIntAdd_group_19: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_635_scaled & simple_obj_ref_634_scaled;
      array_obj_ref_636_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_636_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_636_index_sum_1_req_1;
      array_obj_ref_636_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_636_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : array_obj_ref_642_index_sum_1 
    ApIntAdd_group_20: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_641_scaled & simple_obj_ref_640_scaled;
      array_obj_ref_642_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_642_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_642_index_sum_1_req_1;
      array_obj_ref_642_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_642_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : array_obj_ref_648_index_sum_1 
    ApIntAdd_group_21: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_647_scaled & simple_obj_ref_646_scaled;
      array_obj_ref_648_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_648_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_648_index_sum_1_req_1;
      array_obj_ref_648_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_648_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : array_obj_ref_660_index_sum_1 
    ApIntAdd_group_22: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_659_scaled & simple_obj_ref_658_scaled;
      array_obj_ref_660_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_660_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_660_index_sum_1_req_1;
      array_obj_ref_660_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_660_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : array_obj_ref_666_index_sum_1 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_665_scaled & simple_obj_ref_664_scaled;
      array_obj_ref_666_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_666_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_666_index_sum_1_req_1;
      array_obj_ref_666_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_666_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : array_obj_ref_672_index_sum_1 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_671_scaled & simple_obj_ref_670_scaled;
      array_obj_ref_672_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_672_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_672_index_sum_1_req_1;
      array_obj_ref_672_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_672_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : array_obj_ref_678_index_sum_1 
    ApIntAdd_group_25: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_677_scaled & simple_obj_ref_676_scaled;
      array_obj_ref_678_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_678_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_678_index_sum_1_req_1;
      array_obj_ref_678_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_678_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : array_obj_ref_684_index_sum_1 
    ApIntAdd_group_26: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_683_scaled & simple_obj_ref_682_scaled;
      array_obj_ref_684_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_684_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_684_index_sum_1_req_1;
      array_obj_ref_684_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_684_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : array_obj_ref_690_index_sum_1 
    ApIntAdd_group_27: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_689_scaled & simple_obj_ref_688_scaled;
      array_obj_ref_690_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_690_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_690_index_sum_1_req_1;
      array_obj_ref_690_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_690_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : array_obj_ref_696_index_sum_1 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_695_scaled & simple_obj_ref_694_scaled;
      array_obj_ref_696_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_696_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_696_index_sum_1_req_1;
      array_obj_ref_696_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_696_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_702_index_sum_1 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_701_scaled & simple_obj_ref_700_scaled;
      array_obj_ref_702_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_702_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_702_index_sum_1_req_1;
      array_obj_ref_702_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_702_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_708_index_sum_1 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_707_scaled & simple_obj_ref_706_scaled;
      array_obj_ref_708_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_708_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_708_index_sum_1_req_1;
      array_obj_ref_708_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_708_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_714_index_sum_1 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_713_scaled & simple_obj_ref_712_scaled;
      array_obj_ref_714_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_714_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_714_index_sum_1_req_1;
      array_obj_ref_714_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_714_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_872_index_sum_1 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_871_scaled & simple_obj_ref_870_scaled;
      array_obj_ref_872_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_872_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_872_index_sum_1_req_1;
      array_obj_ref_872_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_872_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : array_obj_ref_884_index_sum_1 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_883_scaled & simple_obj_ref_882_scaled;
      array_obj_ref_884_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_884_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_884_index_sum_1_req_1;
      array_obj_ref_884_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_884_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : array_obj_ref_896_index_sum_1 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_895_scaled & simple_obj_ref_894_scaled;
      array_obj_ref_896_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_896_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_896_index_sum_1_req_1;
      array_obj_ref_896_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_896_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_902_index_sum_1 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_901_scaled & simple_obj_ref_900_scaled;
      array_obj_ref_902_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_902_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_902_index_sum_1_req_1;
      array_obj_ref_902_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_902_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_908_index_sum_1 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_907_scaled & simple_obj_ref_906_scaled;
      array_obj_ref_908_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_908_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_908_index_sum_1_req_1;
      array_obj_ref_908_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_908_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : array_obj_ref_914_index_sum_1 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_913_scaled & simple_obj_ref_912_scaled;
      array_obj_ref_914_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_914_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_914_index_sum_1_req_1;
      array_obj_ref_914_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_914_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : array_obj_ref_926_index_sum_1 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_925_scaled & simple_obj_ref_924_scaled;
      array_obj_ref_926_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_926_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_926_index_sum_1_req_1;
      array_obj_ref_926_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_926_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : array_obj_ref_932_index_sum_1 
    ApIntAdd_group_39: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_931_scaled & simple_obj_ref_930_scaled;
      array_obj_ref_932_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_932_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_932_index_sum_1_req_1;
      array_obj_ref_932_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_932_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : array_obj_ref_938_index_sum_1 
    ApIntAdd_group_40: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_937_scaled & simple_obj_ref_936_scaled;
      array_obj_ref_938_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_938_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_938_index_sum_1_req_1;
      array_obj_ref_938_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_938_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : array_obj_ref_944_index_sum_1 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_943_scaled & simple_obj_ref_942_scaled;
      array_obj_ref_944_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_944_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_944_index_sum_1_req_1;
      array_obj_ref_944_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_944_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : array_obj_ref_950_index_sum_1 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_949_scaled & simple_obj_ref_948_scaled;
      array_obj_ref_950_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_950_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_950_index_sum_1_req_1;
      array_obj_ref_950_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_950_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : array_obj_ref_956_index_sum_1 
    ApIntAdd_group_43: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_955_scaled & simple_obj_ref_954_scaled;
      array_obj_ref_956_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_956_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_956_index_sum_1_req_1;
      array_obj_ref_956_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_956_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : array_obj_ref_962_index_sum_1 
    ApIntAdd_group_44: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_961_scaled & simple_obj_ref_960_scaled;
      array_obj_ref_962_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_962_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_962_index_sum_1_req_1;
      array_obj_ref_962_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_962_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : array_obj_ref_968_index_sum_1 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_967_scaled & simple_obj_ref_966_scaled;
      array_obj_ref_968_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_968_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_968_index_sum_1_req_1;
      array_obj_ref_968_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_968_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : array_obj_ref_974_index_sum_1 
    ApIntAdd_group_46: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_973_scaled & simple_obj_ref_972_scaled;
      array_obj_ref_974_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_974_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_974_index_sum_1_req_1;
      array_obj_ref_974_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_974_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : array_obj_ref_980_index_sum_1 
    ApIntAdd_group_47: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_979_scaled & simple_obj_ref_978_scaled;
      array_obj_ref_980_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_980_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_980_index_sum_1_req_1;
      array_obj_ref_980_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_980_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : array_obj_ref_998_index_sum_1 
    ApIntAdd_group_48: Block -- 
      signal data_in: std_logic_vector(17 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_997_scaled & simple_obj_ref_996_scaled;
      array_obj_ref_998_index_partial_sum_1 <= data_out(8 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= array_obj_ref_998_index_sum_1_req_0;
      reqR(0) <= array_obj_ref_998_index_sum_1_req_1;
      array_obj_ref_998_index_sum_1_ack_0 <= ackL(0); 
      array_obj_ref_998_index_sum_1_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 9, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_1005_inst 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp266_988;
      tmp270_1006 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_1005_inst_req_0;
      reqR(0) <= binary_1005_inst_req_1;
      binary_1005_inst_ack_0 <= ackL(0); 
      binary_1005_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_1017_inst 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp266_988;
      tmp272_1018 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_1017_inst_req_0;
      reqR(0) <= binary_1017_inst_req_1;
      binary_1017_inst_ack_0 <= ackL(0); 
      binary_1017_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_1854_inst binary_1799_inst binary_1794_inst binary_1678_inst binary_1839_inst binary_1834_inst binary_1769_inst binary_1809_inst binary_1814_inst binary_1623_inst binary_1618_inst binary_1754_inst binary_1658_inst binary_1774_inst binary_1849_inst binary_1759_inst binary_1638_inst binary_1633_inst binary_1714_inst binary_1719_inst binary_1729_inst binary_1673_inst binary_1734_inst binary_1663_inst binary_1138_inst binary_1143_inst binary_1153_inst binary_1158_inst binary_1194_inst binary_1199_inst binary_1209_inst binary_1214_inst binary_1250_inst binary_1255_inst binary_1265_inst binary_1270_inst binary_1306_inst binary_1311_inst binary_1321_inst binary_1326_inst binary_1362_inst binary_1367_inst binary_1377_inst binary_1382_inst binary_1402_inst binary_1407_inst binary_1417_inst binary_1422_inst binary_1442_inst binary_1447_inst binary_1457_inst binary_1462_inst binary_1482_inst binary_1487_inst binary_1497_inst binary_1502_inst binary_1538_inst binary_1543_inst binary_1553_inst binary_1558_inst binary_1578_inst binary_1583_inst binary_1593_inst binary_1598_inst 
    ApFloatMul_group_51: Block -- 
      signal data_in: std_logic_vector(4095 downto 0);
      signal data_out: std_logic_vector(2047 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 63 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 63 downto 0);
      signal guard_vector : std_logic_vector( 63 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_130_1710 & iNsTr_46_1302 & iNsTr_128_1702 & iNsTr_32_1238 & iNsTr_127_1698 & iNsTr_31_1234 & iNsTr_94_1534 & iNsTr_46_1302 & iNsTr_128_1702 & iNsTr_44_1294 & iNsTr_127_1698 & iNsTr_43_1290 & iNsTr_129_1706 & iNsTr_21_1186 & iNsTr_129_1706 & iNsTr_33_1242 & iNsTr_130_1710 & iNsTr_34_1246 & iNsTr_92_1526 & iNsTr_32_1238 & iNsTr_91_1522 & iNsTr_31_1234 & iNsTr_127_1698 & iNsTr_19_1178 & iNsTr_91_1522 & iNsTr_43_1290 & iNsTr_130_1710 & iNsTr_22_1190 & iNsTr_129_1706 & iNsTr_45_1298 & iNsTr_128_1702 & iNsTr_20_1182 & iNsTr_94_1534 & iNsTr_34_1246 & iNsTr_93_1530 & iNsTr_33_1242 & iNsTr_127_1698 & iNsTr_4_1110 & iNsTr_128_1702 & iNsTr_6_1118 & iNsTr_129_1706 & iNsTr_8_1126 & iNsTr_93_1530 & iNsTr_45_1298 & iNsTr_130_1710 & iNsTr_10_1134 & iNsTr_92_1526 & iNsTr_44_1294 & iNsTr_3_1106 & iNsTr_4_1110 & iNsTr_5_1114 & iNsTr_6_1118 & iNsTr_7_1122 & iNsTr_8_1126 & iNsTr_9_1130 & iNsTr_10_1134 & iNsTr_3_1106 & iNsTr_19_1178 & iNsTr_5_1114 & iNsTr_20_1182 & iNsTr_7_1122 & iNsTr_21_1186 & iNsTr_9_1130 & iNsTr_22_1190 & iNsTr_3_1106 & iNsTr_31_1234 & iNsTr_5_1114 & iNsTr_32_1238 & iNsTr_7_1122 & iNsTr_33_1242 & iNsTr_9_1130 & iNsTr_34_1246 & iNsTr_3_1106 & iNsTr_43_1290 & iNsTr_5_1114 & iNsTr_44_1294 & iNsTr_7_1122 & iNsTr_45_1298 & iNsTr_9_1130 & iNsTr_46_1302 & iNsTr_55_1346 & iNsTr_4_1110 & iNsTr_56_1350 & iNsTr_6_1118 & iNsTr_57_1354 & iNsTr_8_1126 & iNsTr_58_1358 & iNsTr_10_1134 & iNsTr_55_1346 & iNsTr_19_1178 & iNsTr_56_1350 & iNsTr_20_1182 & iNsTr_57_1354 & iNsTr_21_1186 & iNsTr_58_1358 & iNsTr_22_1190 & iNsTr_55_1346 & iNsTr_31_1234 & iNsTr_56_1350 & iNsTr_32_1238 & iNsTr_57_1354 & iNsTr_33_1242 & iNsTr_58_1358 & iNsTr_34_1246 & iNsTr_55_1346 & iNsTr_43_1290 & iNsTr_56_1350 & iNsTr_44_1294 & iNsTr_57_1354 & iNsTr_45_1298 & iNsTr_58_1358 & iNsTr_46_1302 & iNsTr_91_1522 & iNsTr_4_1110 & iNsTr_92_1526 & iNsTr_6_1118 & iNsTr_93_1530 & iNsTr_8_1126 & iNsTr_94_1534 & iNsTr_10_1134 & iNsTr_91_1522 & iNsTr_19_1178 & iNsTr_92_1526 & iNsTr_20_1182 & iNsTr_93_1530 & iNsTr_21_1186 & iNsTr_94_1534 & iNsTr_22_1190;
      iNsTr_159_1855 <= data_out(2047 downto 2016);
      iNsTr_148_1800 <= data_out(2015 downto 1984);
      iNsTr_147_1795 <= data_out(1983 downto 1952);
      iNsTr_123_1679 <= data_out(1951 downto 1920);
      iNsTr_156_1840 <= data_out(1919 downto 1888);
      iNsTr_155_1835 <= data_out(1887 downto 1856);
      iNsTr_142_1770 <= data_out(1855 downto 1824);
      iNsTr_150_1810 <= data_out(1823 downto 1792);
      iNsTr_151_1815 <= data_out(1791 downto 1760);
      iNsTr_112_1624 <= data_out(1759 downto 1728);
      iNsTr_111_1619 <= data_out(1727 downto 1696);
      iNsTr_139_1755 <= data_out(1695 downto 1664);
      iNsTr_119_1659 <= data_out(1663 downto 1632);
      iNsTr_143_1775 <= data_out(1631 downto 1600);
      iNsTr_158_1850 <= data_out(1599 downto 1568);
      iNsTr_140_1760 <= data_out(1567 downto 1536);
      iNsTr_115_1639 <= data_out(1535 downto 1504);
      iNsTr_114_1634 <= data_out(1503 downto 1472);
      iNsTr_131_1715 <= data_out(1471 downto 1440);
      iNsTr_132_1720 <= data_out(1439 downto 1408);
      iNsTr_134_1730 <= data_out(1407 downto 1376);
      iNsTr_122_1674 <= data_out(1375 downto 1344);
      iNsTr_135_1735 <= data_out(1343 downto 1312);
      iNsTr_120_1664 <= data_out(1311 downto 1280);
      iNsTr_11_1139 <= data_out(1279 downto 1248);
      iNsTr_12_1144 <= data_out(1247 downto 1216);
      iNsTr_14_1154 <= data_out(1215 downto 1184);
      iNsTr_15_1159 <= data_out(1183 downto 1152);
      iNsTr_23_1195 <= data_out(1151 downto 1120);
      iNsTr_24_1200 <= data_out(1119 downto 1088);
      iNsTr_26_1210 <= data_out(1087 downto 1056);
      iNsTr_27_1215 <= data_out(1055 downto 1024);
      iNsTr_35_1251 <= data_out(1023 downto 992);
      iNsTr_36_1256 <= data_out(991 downto 960);
      iNsTr_38_1266 <= data_out(959 downto 928);
      iNsTr_39_1271 <= data_out(927 downto 896);
      iNsTr_47_1307 <= data_out(895 downto 864);
      iNsTr_48_1312 <= data_out(863 downto 832);
      iNsTr_50_1322 <= data_out(831 downto 800);
      iNsTr_51_1327 <= data_out(799 downto 768);
      iNsTr_59_1363 <= data_out(767 downto 736);
      iNsTr_60_1368 <= data_out(735 downto 704);
      iNsTr_62_1378 <= data_out(703 downto 672);
      iNsTr_63_1383 <= data_out(671 downto 640);
      iNsTr_67_1403 <= data_out(639 downto 608);
      iNsTr_68_1408 <= data_out(607 downto 576);
      iNsTr_70_1418 <= data_out(575 downto 544);
      iNsTr_71_1423 <= data_out(543 downto 512);
      iNsTr_75_1443 <= data_out(511 downto 480);
      iNsTr_76_1448 <= data_out(479 downto 448);
      iNsTr_78_1458 <= data_out(447 downto 416);
      iNsTr_79_1463 <= data_out(415 downto 384);
      iNsTr_83_1483 <= data_out(383 downto 352);
      iNsTr_84_1488 <= data_out(351 downto 320);
      iNsTr_86_1498 <= data_out(319 downto 288);
      iNsTr_87_1503 <= data_out(287 downto 256);
      iNsTr_95_1539 <= data_out(255 downto 224);
      iNsTr_96_1544 <= data_out(223 downto 192);
      iNsTr_98_1554 <= data_out(191 downto 160);
      iNsTr_99_1559 <= data_out(159 downto 128);
      iNsTr_103_1579 <= data_out(127 downto 96);
      iNsTr_104_1584 <= data_out(95 downto 64);
      iNsTr_106_1594 <= data_out(63 downto 32);
      iNsTr_107_1599 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      guard_vector(40)  <=  '1';
      guard_vector(41)  <=  '1';
      guard_vector(42)  <=  '1';
      guard_vector(43)  <=  '1';
      guard_vector(44)  <=  '1';
      guard_vector(45)  <=  '1';
      guard_vector(46)  <=  '1';
      guard_vector(47)  <=  '1';
      guard_vector(48)  <=  '1';
      guard_vector(49)  <=  '1';
      guard_vector(50)  <=  '1';
      guard_vector(51)  <=  '1';
      guard_vector(52)  <=  '1';
      guard_vector(53)  <=  '1';
      guard_vector(54)  <=  '1';
      guard_vector(55)  <=  '1';
      guard_vector(56)  <=  '1';
      guard_vector(57)  <=  '1';
      guard_vector(58)  <=  '1';
      guard_vector(59)  <=  '1';
      guard_vector(60)  <=  '1';
      guard_vector(61)  <=  '1';
      guard_vector(62)  <=  '1';
      guard_vector(63)  <=  '1';
      reqL_unguarded(63) <= binary_1854_inst_req_0;
      reqL_unguarded(62) <= binary_1799_inst_req_0;
      reqL_unguarded(61) <= binary_1794_inst_req_0;
      reqL_unguarded(60) <= binary_1678_inst_req_0;
      reqL_unguarded(59) <= binary_1839_inst_req_0;
      reqL_unguarded(58) <= binary_1834_inst_req_0;
      reqL_unguarded(57) <= binary_1769_inst_req_0;
      reqL_unguarded(56) <= binary_1809_inst_req_0;
      reqL_unguarded(55) <= binary_1814_inst_req_0;
      reqL_unguarded(54) <= binary_1623_inst_req_0;
      reqL_unguarded(53) <= binary_1618_inst_req_0;
      reqL_unguarded(52) <= binary_1754_inst_req_0;
      reqL_unguarded(51) <= binary_1658_inst_req_0;
      reqL_unguarded(50) <= binary_1774_inst_req_0;
      reqL_unguarded(49) <= binary_1849_inst_req_0;
      reqL_unguarded(48) <= binary_1759_inst_req_0;
      reqL_unguarded(47) <= binary_1638_inst_req_0;
      reqL_unguarded(46) <= binary_1633_inst_req_0;
      reqL_unguarded(45) <= binary_1714_inst_req_0;
      reqL_unguarded(44) <= binary_1719_inst_req_0;
      reqL_unguarded(43) <= binary_1729_inst_req_0;
      reqL_unguarded(42) <= binary_1673_inst_req_0;
      reqL_unguarded(41) <= binary_1734_inst_req_0;
      reqL_unguarded(40) <= binary_1663_inst_req_0;
      reqL_unguarded(39) <= binary_1138_inst_req_0;
      reqL_unguarded(38) <= binary_1143_inst_req_0;
      reqL_unguarded(37) <= binary_1153_inst_req_0;
      reqL_unguarded(36) <= binary_1158_inst_req_0;
      reqL_unguarded(35) <= binary_1194_inst_req_0;
      reqL_unguarded(34) <= binary_1199_inst_req_0;
      reqL_unguarded(33) <= binary_1209_inst_req_0;
      reqL_unguarded(32) <= binary_1214_inst_req_0;
      reqL_unguarded(31) <= binary_1250_inst_req_0;
      reqL_unguarded(30) <= binary_1255_inst_req_0;
      reqL_unguarded(29) <= binary_1265_inst_req_0;
      reqL_unguarded(28) <= binary_1270_inst_req_0;
      reqL_unguarded(27) <= binary_1306_inst_req_0;
      reqL_unguarded(26) <= binary_1311_inst_req_0;
      reqL_unguarded(25) <= binary_1321_inst_req_0;
      reqL_unguarded(24) <= binary_1326_inst_req_0;
      reqL_unguarded(23) <= binary_1362_inst_req_0;
      reqL_unguarded(22) <= binary_1367_inst_req_0;
      reqL_unguarded(21) <= binary_1377_inst_req_0;
      reqL_unguarded(20) <= binary_1382_inst_req_0;
      reqL_unguarded(19) <= binary_1402_inst_req_0;
      reqL_unguarded(18) <= binary_1407_inst_req_0;
      reqL_unguarded(17) <= binary_1417_inst_req_0;
      reqL_unguarded(16) <= binary_1422_inst_req_0;
      reqL_unguarded(15) <= binary_1442_inst_req_0;
      reqL_unguarded(14) <= binary_1447_inst_req_0;
      reqL_unguarded(13) <= binary_1457_inst_req_0;
      reqL_unguarded(12) <= binary_1462_inst_req_0;
      reqL_unguarded(11) <= binary_1482_inst_req_0;
      reqL_unguarded(10) <= binary_1487_inst_req_0;
      reqL_unguarded(9) <= binary_1497_inst_req_0;
      reqL_unguarded(8) <= binary_1502_inst_req_0;
      reqL_unguarded(7) <= binary_1538_inst_req_0;
      reqL_unguarded(6) <= binary_1543_inst_req_0;
      reqL_unguarded(5) <= binary_1553_inst_req_0;
      reqL_unguarded(4) <= binary_1558_inst_req_0;
      reqL_unguarded(3) <= binary_1578_inst_req_0;
      reqL_unguarded(2) <= binary_1583_inst_req_0;
      reqL_unguarded(1) <= binary_1593_inst_req_0;
      reqL_unguarded(0) <= binary_1598_inst_req_0;
      binary_1854_inst_ack_0 <= ackL_unguarded(63);
      binary_1799_inst_ack_0 <= ackL_unguarded(62);
      binary_1794_inst_ack_0 <= ackL_unguarded(61);
      binary_1678_inst_ack_0 <= ackL_unguarded(60);
      binary_1839_inst_ack_0 <= ackL_unguarded(59);
      binary_1834_inst_ack_0 <= ackL_unguarded(58);
      binary_1769_inst_ack_0 <= ackL_unguarded(57);
      binary_1809_inst_ack_0 <= ackL_unguarded(56);
      binary_1814_inst_ack_0 <= ackL_unguarded(55);
      binary_1623_inst_ack_0 <= ackL_unguarded(54);
      binary_1618_inst_ack_0 <= ackL_unguarded(53);
      binary_1754_inst_ack_0 <= ackL_unguarded(52);
      binary_1658_inst_ack_0 <= ackL_unguarded(51);
      binary_1774_inst_ack_0 <= ackL_unguarded(50);
      binary_1849_inst_ack_0 <= ackL_unguarded(49);
      binary_1759_inst_ack_0 <= ackL_unguarded(48);
      binary_1638_inst_ack_0 <= ackL_unguarded(47);
      binary_1633_inst_ack_0 <= ackL_unguarded(46);
      binary_1714_inst_ack_0 <= ackL_unguarded(45);
      binary_1719_inst_ack_0 <= ackL_unguarded(44);
      binary_1729_inst_ack_0 <= ackL_unguarded(43);
      binary_1673_inst_ack_0 <= ackL_unguarded(42);
      binary_1734_inst_ack_0 <= ackL_unguarded(41);
      binary_1663_inst_ack_0 <= ackL_unguarded(40);
      binary_1138_inst_ack_0 <= ackL_unguarded(39);
      binary_1143_inst_ack_0 <= ackL_unguarded(38);
      binary_1153_inst_ack_0 <= ackL_unguarded(37);
      binary_1158_inst_ack_0 <= ackL_unguarded(36);
      binary_1194_inst_ack_0 <= ackL_unguarded(35);
      binary_1199_inst_ack_0 <= ackL_unguarded(34);
      binary_1209_inst_ack_0 <= ackL_unguarded(33);
      binary_1214_inst_ack_0 <= ackL_unguarded(32);
      binary_1250_inst_ack_0 <= ackL_unguarded(31);
      binary_1255_inst_ack_0 <= ackL_unguarded(30);
      binary_1265_inst_ack_0 <= ackL_unguarded(29);
      binary_1270_inst_ack_0 <= ackL_unguarded(28);
      binary_1306_inst_ack_0 <= ackL_unguarded(27);
      binary_1311_inst_ack_0 <= ackL_unguarded(26);
      binary_1321_inst_ack_0 <= ackL_unguarded(25);
      binary_1326_inst_ack_0 <= ackL_unguarded(24);
      binary_1362_inst_ack_0 <= ackL_unguarded(23);
      binary_1367_inst_ack_0 <= ackL_unguarded(22);
      binary_1377_inst_ack_0 <= ackL_unguarded(21);
      binary_1382_inst_ack_0 <= ackL_unguarded(20);
      binary_1402_inst_ack_0 <= ackL_unguarded(19);
      binary_1407_inst_ack_0 <= ackL_unguarded(18);
      binary_1417_inst_ack_0 <= ackL_unguarded(17);
      binary_1422_inst_ack_0 <= ackL_unguarded(16);
      binary_1442_inst_ack_0 <= ackL_unguarded(15);
      binary_1447_inst_ack_0 <= ackL_unguarded(14);
      binary_1457_inst_ack_0 <= ackL_unguarded(13);
      binary_1462_inst_ack_0 <= ackL_unguarded(12);
      binary_1482_inst_ack_0 <= ackL_unguarded(11);
      binary_1487_inst_ack_0 <= ackL_unguarded(10);
      binary_1497_inst_ack_0 <= ackL_unguarded(9);
      binary_1502_inst_ack_0 <= ackL_unguarded(8);
      binary_1538_inst_ack_0 <= ackL_unguarded(7);
      binary_1543_inst_ack_0 <= ackL_unguarded(6);
      binary_1553_inst_ack_0 <= ackL_unguarded(5);
      binary_1558_inst_ack_0 <= ackL_unguarded(4);
      binary_1578_inst_ack_0 <= ackL_unguarded(3);
      binary_1583_inst_ack_0 <= ackL_unguarded(2);
      binary_1593_inst_ack_0 <= ackL_unguarded(1);
      binary_1598_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(63) <= binary_1854_inst_req_1;
      reqR_unguarded(62) <= binary_1799_inst_req_1;
      reqR_unguarded(61) <= binary_1794_inst_req_1;
      reqR_unguarded(60) <= binary_1678_inst_req_1;
      reqR_unguarded(59) <= binary_1839_inst_req_1;
      reqR_unguarded(58) <= binary_1834_inst_req_1;
      reqR_unguarded(57) <= binary_1769_inst_req_1;
      reqR_unguarded(56) <= binary_1809_inst_req_1;
      reqR_unguarded(55) <= binary_1814_inst_req_1;
      reqR_unguarded(54) <= binary_1623_inst_req_1;
      reqR_unguarded(53) <= binary_1618_inst_req_1;
      reqR_unguarded(52) <= binary_1754_inst_req_1;
      reqR_unguarded(51) <= binary_1658_inst_req_1;
      reqR_unguarded(50) <= binary_1774_inst_req_1;
      reqR_unguarded(49) <= binary_1849_inst_req_1;
      reqR_unguarded(48) <= binary_1759_inst_req_1;
      reqR_unguarded(47) <= binary_1638_inst_req_1;
      reqR_unguarded(46) <= binary_1633_inst_req_1;
      reqR_unguarded(45) <= binary_1714_inst_req_1;
      reqR_unguarded(44) <= binary_1719_inst_req_1;
      reqR_unguarded(43) <= binary_1729_inst_req_1;
      reqR_unguarded(42) <= binary_1673_inst_req_1;
      reqR_unguarded(41) <= binary_1734_inst_req_1;
      reqR_unguarded(40) <= binary_1663_inst_req_1;
      reqR_unguarded(39) <= binary_1138_inst_req_1;
      reqR_unguarded(38) <= binary_1143_inst_req_1;
      reqR_unguarded(37) <= binary_1153_inst_req_1;
      reqR_unguarded(36) <= binary_1158_inst_req_1;
      reqR_unguarded(35) <= binary_1194_inst_req_1;
      reqR_unguarded(34) <= binary_1199_inst_req_1;
      reqR_unguarded(33) <= binary_1209_inst_req_1;
      reqR_unguarded(32) <= binary_1214_inst_req_1;
      reqR_unguarded(31) <= binary_1250_inst_req_1;
      reqR_unguarded(30) <= binary_1255_inst_req_1;
      reqR_unguarded(29) <= binary_1265_inst_req_1;
      reqR_unguarded(28) <= binary_1270_inst_req_1;
      reqR_unguarded(27) <= binary_1306_inst_req_1;
      reqR_unguarded(26) <= binary_1311_inst_req_1;
      reqR_unguarded(25) <= binary_1321_inst_req_1;
      reqR_unguarded(24) <= binary_1326_inst_req_1;
      reqR_unguarded(23) <= binary_1362_inst_req_1;
      reqR_unguarded(22) <= binary_1367_inst_req_1;
      reqR_unguarded(21) <= binary_1377_inst_req_1;
      reqR_unguarded(20) <= binary_1382_inst_req_1;
      reqR_unguarded(19) <= binary_1402_inst_req_1;
      reqR_unguarded(18) <= binary_1407_inst_req_1;
      reqR_unguarded(17) <= binary_1417_inst_req_1;
      reqR_unguarded(16) <= binary_1422_inst_req_1;
      reqR_unguarded(15) <= binary_1442_inst_req_1;
      reqR_unguarded(14) <= binary_1447_inst_req_1;
      reqR_unguarded(13) <= binary_1457_inst_req_1;
      reqR_unguarded(12) <= binary_1462_inst_req_1;
      reqR_unguarded(11) <= binary_1482_inst_req_1;
      reqR_unguarded(10) <= binary_1487_inst_req_1;
      reqR_unguarded(9) <= binary_1497_inst_req_1;
      reqR_unguarded(8) <= binary_1502_inst_req_1;
      reqR_unguarded(7) <= binary_1538_inst_req_1;
      reqR_unguarded(6) <= binary_1543_inst_req_1;
      reqR_unguarded(5) <= binary_1553_inst_req_1;
      reqR_unguarded(4) <= binary_1558_inst_req_1;
      reqR_unguarded(3) <= binary_1578_inst_req_1;
      reqR_unguarded(2) <= binary_1583_inst_req_1;
      reqR_unguarded(1) <= binary_1593_inst_req_1;
      reqR_unguarded(0) <= binary_1598_inst_req_1;
      binary_1854_inst_ack_1 <= ackR_unguarded(63);
      binary_1799_inst_ack_1 <= ackR_unguarded(62);
      binary_1794_inst_ack_1 <= ackR_unguarded(61);
      binary_1678_inst_ack_1 <= ackR_unguarded(60);
      binary_1839_inst_ack_1 <= ackR_unguarded(59);
      binary_1834_inst_ack_1 <= ackR_unguarded(58);
      binary_1769_inst_ack_1 <= ackR_unguarded(57);
      binary_1809_inst_ack_1 <= ackR_unguarded(56);
      binary_1814_inst_ack_1 <= ackR_unguarded(55);
      binary_1623_inst_ack_1 <= ackR_unguarded(54);
      binary_1618_inst_ack_1 <= ackR_unguarded(53);
      binary_1754_inst_ack_1 <= ackR_unguarded(52);
      binary_1658_inst_ack_1 <= ackR_unguarded(51);
      binary_1774_inst_ack_1 <= ackR_unguarded(50);
      binary_1849_inst_ack_1 <= ackR_unguarded(49);
      binary_1759_inst_ack_1 <= ackR_unguarded(48);
      binary_1638_inst_ack_1 <= ackR_unguarded(47);
      binary_1633_inst_ack_1 <= ackR_unguarded(46);
      binary_1714_inst_ack_1 <= ackR_unguarded(45);
      binary_1719_inst_ack_1 <= ackR_unguarded(44);
      binary_1729_inst_ack_1 <= ackR_unguarded(43);
      binary_1673_inst_ack_1 <= ackR_unguarded(42);
      binary_1734_inst_ack_1 <= ackR_unguarded(41);
      binary_1663_inst_ack_1 <= ackR_unguarded(40);
      binary_1138_inst_ack_1 <= ackR_unguarded(39);
      binary_1143_inst_ack_1 <= ackR_unguarded(38);
      binary_1153_inst_ack_1 <= ackR_unguarded(37);
      binary_1158_inst_ack_1 <= ackR_unguarded(36);
      binary_1194_inst_ack_1 <= ackR_unguarded(35);
      binary_1199_inst_ack_1 <= ackR_unguarded(34);
      binary_1209_inst_ack_1 <= ackR_unguarded(33);
      binary_1214_inst_ack_1 <= ackR_unguarded(32);
      binary_1250_inst_ack_1 <= ackR_unguarded(31);
      binary_1255_inst_ack_1 <= ackR_unguarded(30);
      binary_1265_inst_ack_1 <= ackR_unguarded(29);
      binary_1270_inst_ack_1 <= ackR_unguarded(28);
      binary_1306_inst_ack_1 <= ackR_unguarded(27);
      binary_1311_inst_ack_1 <= ackR_unguarded(26);
      binary_1321_inst_ack_1 <= ackR_unguarded(25);
      binary_1326_inst_ack_1 <= ackR_unguarded(24);
      binary_1362_inst_ack_1 <= ackR_unguarded(23);
      binary_1367_inst_ack_1 <= ackR_unguarded(22);
      binary_1377_inst_ack_1 <= ackR_unguarded(21);
      binary_1382_inst_ack_1 <= ackR_unguarded(20);
      binary_1402_inst_ack_1 <= ackR_unguarded(19);
      binary_1407_inst_ack_1 <= ackR_unguarded(18);
      binary_1417_inst_ack_1 <= ackR_unguarded(17);
      binary_1422_inst_ack_1 <= ackR_unguarded(16);
      binary_1442_inst_ack_1 <= ackR_unguarded(15);
      binary_1447_inst_ack_1 <= ackR_unguarded(14);
      binary_1457_inst_ack_1 <= ackR_unguarded(13);
      binary_1462_inst_ack_1 <= ackR_unguarded(12);
      binary_1482_inst_ack_1 <= ackR_unguarded(11);
      binary_1487_inst_ack_1 <= ackR_unguarded(10);
      binary_1497_inst_ack_1 <= ackR_unguarded(9);
      binary_1502_inst_ack_1 <= ackR_unguarded(8);
      binary_1538_inst_ack_1 <= ackR_unguarded(7);
      binary_1543_inst_ack_1 <= ackR_unguarded(6);
      binary_1553_inst_ack_1 <= ackR_unguarded(5);
      binary_1558_inst_ack_1 <= ackR_unguarded(4);
      binary_1578_inst_ack_1 <= ackR_unguarded(3);
      binary_1583_inst_ack_1 <= ackR_unguarded(2);
      binary_1593_inst_ack_1 <= ackR_unguarded(1);
      binary_1598_inst_ack_1 <= ackR_unguarded(0);
      gI0: GuardInterface generic map(nreqs => 64) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 64) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          operator_id => "ApFloatMul",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 64 -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_1844_inst binary_1764_inst binary_1608_inst binary_1789_inst binary_1784_inst binary_1829_inst binary_1859_inst binary_1864_inst binary_1824_inst binary_1693_inst binary_1819_inst binary_1779_inst binary_1869_inst binary_1683_inst binary_1628_inst binary_1643_inst binary_1613_inst binary_1688_inst binary_1648_inst binary_1653_inst binary_1724_inst binary_1739_inst binary_1744_inst binary_1749_inst binary_1668_inst binary_1804_inst binary_1148_inst binary_1163_inst binary_1168_inst binary_1173_inst binary_1204_inst binary_1219_inst binary_1224_inst binary_1229_inst binary_1260_inst binary_1275_inst binary_1280_inst binary_1285_inst binary_1316_inst binary_1331_inst binary_1336_inst binary_1341_inst binary_1372_inst binary_1387_inst binary_1392_inst binary_1397_inst binary_1412_inst binary_1427_inst binary_1432_inst binary_1437_inst binary_1452_inst binary_1467_inst binary_1472_inst binary_1477_inst binary_1492_inst binary_1507_inst binary_1512_inst binary_1517_inst binary_1548_inst binary_1563_inst binary_1568_inst binary_1573_inst binary_1588_inst binary_1603_inst 
    ApFloatAdd_group_52: Block -- 
      signal data_in: std_logic_vector(4095 downto 0);
      signal data_out: std_logic_vector(2047 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 63 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 63 downto 0);
      signal guard_vector : std_logic_vector( 63 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_155_1835 & iNsTr_156_1840 & iNsTr_139_1755 & iNsTr_140_1760 & iNsTr_105_1589 & iNsTr_108_1604 & v31x_x016_764 & iNsTr_145_1785 & iNsTr_141_1765 & iNsTr_144_1780 & v32x_x017_757 & iNsTr_153_1825 & iNsTr_158_1850 & iNsTr_159_1855 & iNsTr_157_1845 & iNsTr_160_1860 & iNsTr_149_1805 & iNsTr_152_1820 & v23x_x014_778 & iNsTr_125_1689 & iNsTr_150_1810 & iNsTr_151_1815 & iNsTr_142_1770 & iNsTr_143_1775 & v33x_x018_750 & iNsTr_161_1865 & iNsTr_122_1674 & iNsTr_123_1679 & iNsTr_111_1619 & iNsTr_112_1624 & iNsTr_114_1634 & iNsTr_115_1639 & v21x_x012_792 & iNsTr_109_1609 & iNsTr_121_1669 & iNsTr_124_1684 & iNsTr_113_1629 & iNsTr_116_1644 & v22x_x013_785 & iNsTr_117_1649 & iNsTr_131_1715 & iNsTr_132_1720 & iNsTr_134_1730 & iNsTr_135_1735 & iNsTr_133_1725 & iNsTr_136_1740 & v30x_x015_771 & iNsTr_137_1745 & iNsTr_119_1659 & iNsTr_120_1664 & iNsTr_147_1795 & iNsTr_148_1800 & iNsTr_11_1139 & iNsTr_12_1144 & iNsTr_14_1154 & iNsTr_15_1159 & iNsTr_13_1149 & iNsTr_16_1164 & v00x_x09_813 & iNsTr_17_1169 & iNsTr_23_1195 & iNsTr_24_1200 & iNsTr_26_1210 & iNsTr_27_1215 & iNsTr_25_1205 & iNsTr_28_1220 & v01x_x08_820 & iNsTr_29_1225 & iNsTr_35_1251 & iNsTr_36_1256 & iNsTr_38_1266 & iNsTr_39_1271 & iNsTr_37_1261 & iNsTr_40_1276 & v02x_x07_827 & iNsTr_41_1281 & iNsTr_47_1307 & iNsTr_48_1312 & iNsTr_50_1322 & iNsTr_51_1327 & iNsTr_49_1317 & iNsTr_52_1332 & v03x_x06_834 & iNsTr_53_1337 & iNsTr_59_1363 & iNsTr_60_1368 & iNsTr_62_1378 & iNsTr_63_1383 & iNsTr_61_1373 & iNsTr_64_1388 & v10x_x05_841 & iNsTr_65_1393 & iNsTr_67_1403 & iNsTr_68_1408 & iNsTr_70_1418 & iNsTr_71_1423 & iNsTr_69_1413 & iNsTr_72_1428 & v11x_x04_848 & iNsTr_73_1433 & iNsTr_75_1443 & iNsTr_76_1448 & iNsTr_78_1458 & iNsTr_79_1463 & iNsTr_77_1453 & iNsTr_80_1468 & v12x_x03_855 & iNsTr_81_1473 & iNsTr_83_1483 & iNsTr_84_1488 & iNsTr_86_1498 & iNsTr_87_1503 & iNsTr_85_1493 & iNsTr_88_1508 & v13x_x010_806 & iNsTr_89_1513 & iNsTr_95_1539 & iNsTr_96_1544 & iNsTr_98_1554 & iNsTr_99_1559 & iNsTr_97_1549 & iNsTr_100_1564 & v20x_x011_799 & iNsTr_101_1569 & iNsTr_103_1579 & iNsTr_104_1584 & iNsTr_106_1594 & iNsTr_107_1599;
      iNsTr_157_1845 <= data_out(2047 downto 2016);
      iNsTr_141_1765 <= data_out(2015 downto 1984);
      iNsTr_109_1609 <= data_out(1983 downto 1952);
      iNsTr_146_1790 <= data_out(1951 downto 1920);
      iNsTr_145_1785 <= data_out(1919 downto 1888);
      iNsTr_154_1830 <= data_out(1887 downto 1856);
      iNsTr_160_1860 <= data_out(1855 downto 1824);
      iNsTr_161_1865 <= data_out(1823 downto 1792);
      iNsTr_153_1825 <= data_out(1791 downto 1760);
      iNsTr_126_1694 <= data_out(1759 downto 1728);
      iNsTr_152_1820 <= data_out(1727 downto 1696);
      iNsTr_144_1780 <= data_out(1695 downto 1664);
      iNsTr_162_1870 <= data_out(1663 downto 1632);
      iNsTr_124_1684 <= data_out(1631 downto 1600);
      iNsTr_113_1629 <= data_out(1599 downto 1568);
      iNsTr_116_1644 <= data_out(1567 downto 1536);
      iNsTr_110_1614 <= data_out(1535 downto 1504);
      iNsTr_125_1689 <= data_out(1503 downto 1472);
      iNsTr_117_1649 <= data_out(1471 downto 1440);
      iNsTr_118_1654 <= data_out(1439 downto 1408);
      iNsTr_133_1725 <= data_out(1407 downto 1376);
      iNsTr_136_1740 <= data_out(1375 downto 1344);
      iNsTr_137_1745 <= data_out(1343 downto 1312);
      iNsTr_138_1750 <= data_out(1311 downto 1280);
      iNsTr_121_1669 <= data_out(1279 downto 1248);
      iNsTr_149_1805 <= data_out(1247 downto 1216);
      iNsTr_13_1149 <= data_out(1215 downto 1184);
      iNsTr_16_1164 <= data_out(1183 downto 1152);
      iNsTr_17_1169 <= data_out(1151 downto 1120);
      iNsTr_18_1174 <= data_out(1119 downto 1088);
      iNsTr_25_1205 <= data_out(1087 downto 1056);
      iNsTr_28_1220 <= data_out(1055 downto 1024);
      iNsTr_29_1225 <= data_out(1023 downto 992);
      iNsTr_30_1230 <= data_out(991 downto 960);
      iNsTr_37_1261 <= data_out(959 downto 928);
      iNsTr_40_1276 <= data_out(927 downto 896);
      iNsTr_41_1281 <= data_out(895 downto 864);
      iNsTr_42_1286 <= data_out(863 downto 832);
      iNsTr_49_1317 <= data_out(831 downto 800);
      iNsTr_52_1332 <= data_out(799 downto 768);
      iNsTr_53_1337 <= data_out(767 downto 736);
      iNsTr_54_1342 <= data_out(735 downto 704);
      iNsTr_61_1373 <= data_out(703 downto 672);
      iNsTr_64_1388 <= data_out(671 downto 640);
      iNsTr_65_1393 <= data_out(639 downto 608);
      iNsTr_66_1398 <= data_out(607 downto 576);
      iNsTr_69_1413 <= data_out(575 downto 544);
      iNsTr_72_1428 <= data_out(543 downto 512);
      iNsTr_73_1433 <= data_out(511 downto 480);
      iNsTr_74_1438 <= data_out(479 downto 448);
      iNsTr_77_1453 <= data_out(447 downto 416);
      iNsTr_80_1468 <= data_out(415 downto 384);
      iNsTr_81_1473 <= data_out(383 downto 352);
      iNsTr_82_1478 <= data_out(351 downto 320);
      iNsTr_85_1493 <= data_out(319 downto 288);
      iNsTr_88_1508 <= data_out(287 downto 256);
      iNsTr_89_1513 <= data_out(255 downto 224);
      iNsTr_90_1518 <= data_out(223 downto 192);
      iNsTr_97_1549 <= data_out(191 downto 160);
      iNsTr_100_1564 <= data_out(159 downto 128);
      iNsTr_101_1569 <= data_out(127 downto 96);
      iNsTr_102_1574 <= data_out(95 downto 64);
      iNsTr_105_1589 <= data_out(63 downto 32);
      iNsTr_108_1604 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      guard_vector(40)  <=  '1';
      guard_vector(41)  <=  '1';
      guard_vector(42)  <=  '1';
      guard_vector(43)  <=  '1';
      guard_vector(44)  <=  '1';
      guard_vector(45)  <=  '1';
      guard_vector(46)  <=  '1';
      guard_vector(47)  <=  '1';
      guard_vector(48)  <=  '1';
      guard_vector(49)  <=  '1';
      guard_vector(50)  <=  '1';
      guard_vector(51)  <=  '1';
      guard_vector(52)  <=  '1';
      guard_vector(53)  <=  '1';
      guard_vector(54)  <=  '1';
      guard_vector(55)  <=  '1';
      guard_vector(56)  <=  '1';
      guard_vector(57)  <=  '1';
      guard_vector(58)  <=  '1';
      guard_vector(59)  <=  '1';
      guard_vector(60)  <=  '1';
      guard_vector(61)  <=  '1';
      guard_vector(62)  <=  '1';
      guard_vector(63)  <=  '1';
      reqL_unguarded(63) <= binary_1844_inst_req_0;
      reqL_unguarded(62) <= binary_1764_inst_req_0;
      reqL_unguarded(61) <= binary_1608_inst_req_0;
      reqL_unguarded(60) <= binary_1789_inst_req_0;
      reqL_unguarded(59) <= binary_1784_inst_req_0;
      reqL_unguarded(58) <= binary_1829_inst_req_0;
      reqL_unguarded(57) <= binary_1859_inst_req_0;
      reqL_unguarded(56) <= binary_1864_inst_req_0;
      reqL_unguarded(55) <= binary_1824_inst_req_0;
      reqL_unguarded(54) <= binary_1693_inst_req_0;
      reqL_unguarded(53) <= binary_1819_inst_req_0;
      reqL_unguarded(52) <= binary_1779_inst_req_0;
      reqL_unguarded(51) <= binary_1869_inst_req_0;
      reqL_unguarded(50) <= binary_1683_inst_req_0;
      reqL_unguarded(49) <= binary_1628_inst_req_0;
      reqL_unguarded(48) <= binary_1643_inst_req_0;
      reqL_unguarded(47) <= binary_1613_inst_req_0;
      reqL_unguarded(46) <= binary_1688_inst_req_0;
      reqL_unguarded(45) <= binary_1648_inst_req_0;
      reqL_unguarded(44) <= binary_1653_inst_req_0;
      reqL_unguarded(43) <= binary_1724_inst_req_0;
      reqL_unguarded(42) <= binary_1739_inst_req_0;
      reqL_unguarded(41) <= binary_1744_inst_req_0;
      reqL_unguarded(40) <= binary_1749_inst_req_0;
      reqL_unguarded(39) <= binary_1668_inst_req_0;
      reqL_unguarded(38) <= binary_1804_inst_req_0;
      reqL_unguarded(37) <= binary_1148_inst_req_0;
      reqL_unguarded(36) <= binary_1163_inst_req_0;
      reqL_unguarded(35) <= binary_1168_inst_req_0;
      reqL_unguarded(34) <= binary_1173_inst_req_0;
      reqL_unguarded(33) <= binary_1204_inst_req_0;
      reqL_unguarded(32) <= binary_1219_inst_req_0;
      reqL_unguarded(31) <= binary_1224_inst_req_0;
      reqL_unguarded(30) <= binary_1229_inst_req_0;
      reqL_unguarded(29) <= binary_1260_inst_req_0;
      reqL_unguarded(28) <= binary_1275_inst_req_0;
      reqL_unguarded(27) <= binary_1280_inst_req_0;
      reqL_unguarded(26) <= binary_1285_inst_req_0;
      reqL_unguarded(25) <= binary_1316_inst_req_0;
      reqL_unguarded(24) <= binary_1331_inst_req_0;
      reqL_unguarded(23) <= binary_1336_inst_req_0;
      reqL_unguarded(22) <= binary_1341_inst_req_0;
      reqL_unguarded(21) <= binary_1372_inst_req_0;
      reqL_unguarded(20) <= binary_1387_inst_req_0;
      reqL_unguarded(19) <= binary_1392_inst_req_0;
      reqL_unguarded(18) <= binary_1397_inst_req_0;
      reqL_unguarded(17) <= binary_1412_inst_req_0;
      reqL_unguarded(16) <= binary_1427_inst_req_0;
      reqL_unguarded(15) <= binary_1432_inst_req_0;
      reqL_unguarded(14) <= binary_1437_inst_req_0;
      reqL_unguarded(13) <= binary_1452_inst_req_0;
      reqL_unguarded(12) <= binary_1467_inst_req_0;
      reqL_unguarded(11) <= binary_1472_inst_req_0;
      reqL_unguarded(10) <= binary_1477_inst_req_0;
      reqL_unguarded(9) <= binary_1492_inst_req_0;
      reqL_unguarded(8) <= binary_1507_inst_req_0;
      reqL_unguarded(7) <= binary_1512_inst_req_0;
      reqL_unguarded(6) <= binary_1517_inst_req_0;
      reqL_unguarded(5) <= binary_1548_inst_req_0;
      reqL_unguarded(4) <= binary_1563_inst_req_0;
      reqL_unguarded(3) <= binary_1568_inst_req_0;
      reqL_unguarded(2) <= binary_1573_inst_req_0;
      reqL_unguarded(1) <= binary_1588_inst_req_0;
      reqL_unguarded(0) <= binary_1603_inst_req_0;
      binary_1844_inst_ack_0 <= ackL_unguarded(63);
      binary_1764_inst_ack_0 <= ackL_unguarded(62);
      binary_1608_inst_ack_0 <= ackL_unguarded(61);
      binary_1789_inst_ack_0 <= ackL_unguarded(60);
      binary_1784_inst_ack_0 <= ackL_unguarded(59);
      binary_1829_inst_ack_0 <= ackL_unguarded(58);
      binary_1859_inst_ack_0 <= ackL_unguarded(57);
      binary_1864_inst_ack_0 <= ackL_unguarded(56);
      binary_1824_inst_ack_0 <= ackL_unguarded(55);
      binary_1693_inst_ack_0 <= ackL_unguarded(54);
      binary_1819_inst_ack_0 <= ackL_unguarded(53);
      binary_1779_inst_ack_0 <= ackL_unguarded(52);
      binary_1869_inst_ack_0 <= ackL_unguarded(51);
      binary_1683_inst_ack_0 <= ackL_unguarded(50);
      binary_1628_inst_ack_0 <= ackL_unguarded(49);
      binary_1643_inst_ack_0 <= ackL_unguarded(48);
      binary_1613_inst_ack_0 <= ackL_unguarded(47);
      binary_1688_inst_ack_0 <= ackL_unguarded(46);
      binary_1648_inst_ack_0 <= ackL_unguarded(45);
      binary_1653_inst_ack_0 <= ackL_unguarded(44);
      binary_1724_inst_ack_0 <= ackL_unguarded(43);
      binary_1739_inst_ack_0 <= ackL_unguarded(42);
      binary_1744_inst_ack_0 <= ackL_unguarded(41);
      binary_1749_inst_ack_0 <= ackL_unguarded(40);
      binary_1668_inst_ack_0 <= ackL_unguarded(39);
      binary_1804_inst_ack_0 <= ackL_unguarded(38);
      binary_1148_inst_ack_0 <= ackL_unguarded(37);
      binary_1163_inst_ack_0 <= ackL_unguarded(36);
      binary_1168_inst_ack_0 <= ackL_unguarded(35);
      binary_1173_inst_ack_0 <= ackL_unguarded(34);
      binary_1204_inst_ack_0 <= ackL_unguarded(33);
      binary_1219_inst_ack_0 <= ackL_unguarded(32);
      binary_1224_inst_ack_0 <= ackL_unguarded(31);
      binary_1229_inst_ack_0 <= ackL_unguarded(30);
      binary_1260_inst_ack_0 <= ackL_unguarded(29);
      binary_1275_inst_ack_0 <= ackL_unguarded(28);
      binary_1280_inst_ack_0 <= ackL_unguarded(27);
      binary_1285_inst_ack_0 <= ackL_unguarded(26);
      binary_1316_inst_ack_0 <= ackL_unguarded(25);
      binary_1331_inst_ack_0 <= ackL_unguarded(24);
      binary_1336_inst_ack_0 <= ackL_unguarded(23);
      binary_1341_inst_ack_0 <= ackL_unguarded(22);
      binary_1372_inst_ack_0 <= ackL_unguarded(21);
      binary_1387_inst_ack_0 <= ackL_unguarded(20);
      binary_1392_inst_ack_0 <= ackL_unguarded(19);
      binary_1397_inst_ack_0 <= ackL_unguarded(18);
      binary_1412_inst_ack_0 <= ackL_unguarded(17);
      binary_1427_inst_ack_0 <= ackL_unguarded(16);
      binary_1432_inst_ack_0 <= ackL_unguarded(15);
      binary_1437_inst_ack_0 <= ackL_unguarded(14);
      binary_1452_inst_ack_0 <= ackL_unguarded(13);
      binary_1467_inst_ack_0 <= ackL_unguarded(12);
      binary_1472_inst_ack_0 <= ackL_unguarded(11);
      binary_1477_inst_ack_0 <= ackL_unguarded(10);
      binary_1492_inst_ack_0 <= ackL_unguarded(9);
      binary_1507_inst_ack_0 <= ackL_unguarded(8);
      binary_1512_inst_ack_0 <= ackL_unguarded(7);
      binary_1517_inst_ack_0 <= ackL_unguarded(6);
      binary_1548_inst_ack_0 <= ackL_unguarded(5);
      binary_1563_inst_ack_0 <= ackL_unguarded(4);
      binary_1568_inst_ack_0 <= ackL_unguarded(3);
      binary_1573_inst_ack_0 <= ackL_unguarded(2);
      binary_1588_inst_ack_0 <= ackL_unguarded(1);
      binary_1603_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(63) <= binary_1844_inst_req_1;
      reqR_unguarded(62) <= binary_1764_inst_req_1;
      reqR_unguarded(61) <= binary_1608_inst_req_1;
      reqR_unguarded(60) <= binary_1789_inst_req_1;
      reqR_unguarded(59) <= binary_1784_inst_req_1;
      reqR_unguarded(58) <= binary_1829_inst_req_1;
      reqR_unguarded(57) <= binary_1859_inst_req_1;
      reqR_unguarded(56) <= binary_1864_inst_req_1;
      reqR_unguarded(55) <= binary_1824_inst_req_1;
      reqR_unguarded(54) <= binary_1693_inst_req_1;
      reqR_unguarded(53) <= binary_1819_inst_req_1;
      reqR_unguarded(52) <= binary_1779_inst_req_1;
      reqR_unguarded(51) <= binary_1869_inst_req_1;
      reqR_unguarded(50) <= binary_1683_inst_req_1;
      reqR_unguarded(49) <= binary_1628_inst_req_1;
      reqR_unguarded(48) <= binary_1643_inst_req_1;
      reqR_unguarded(47) <= binary_1613_inst_req_1;
      reqR_unguarded(46) <= binary_1688_inst_req_1;
      reqR_unguarded(45) <= binary_1648_inst_req_1;
      reqR_unguarded(44) <= binary_1653_inst_req_1;
      reqR_unguarded(43) <= binary_1724_inst_req_1;
      reqR_unguarded(42) <= binary_1739_inst_req_1;
      reqR_unguarded(41) <= binary_1744_inst_req_1;
      reqR_unguarded(40) <= binary_1749_inst_req_1;
      reqR_unguarded(39) <= binary_1668_inst_req_1;
      reqR_unguarded(38) <= binary_1804_inst_req_1;
      reqR_unguarded(37) <= binary_1148_inst_req_1;
      reqR_unguarded(36) <= binary_1163_inst_req_1;
      reqR_unguarded(35) <= binary_1168_inst_req_1;
      reqR_unguarded(34) <= binary_1173_inst_req_1;
      reqR_unguarded(33) <= binary_1204_inst_req_1;
      reqR_unguarded(32) <= binary_1219_inst_req_1;
      reqR_unguarded(31) <= binary_1224_inst_req_1;
      reqR_unguarded(30) <= binary_1229_inst_req_1;
      reqR_unguarded(29) <= binary_1260_inst_req_1;
      reqR_unguarded(28) <= binary_1275_inst_req_1;
      reqR_unguarded(27) <= binary_1280_inst_req_1;
      reqR_unguarded(26) <= binary_1285_inst_req_1;
      reqR_unguarded(25) <= binary_1316_inst_req_1;
      reqR_unguarded(24) <= binary_1331_inst_req_1;
      reqR_unguarded(23) <= binary_1336_inst_req_1;
      reqR_unguarded(22) <= binary_1341_inst_req_1;
      reqR_unguarded(21) <= binary_1372_inst_req_1;
      reqR_unguarded(20) <= binary_1387_inst_req_1;
      reqR_unguarded(19) <= binary_1392_inst_req_1;
      reqR_unguarded(18) <= binary_1397_inst_req_1;
      reqR_unguarded(17) <= binary_1412_inst_req_1;
      reqR_unguarded(16) <= binary_1427_inst_req_1;
      reqR_unguarded(15) <= binary_1432_inst_req_1;
      reqR_unguarded(14) <= binary_1437_inst_req_1;
      reqR_unguarded(13) <= binary_1452_inst_req_1;
      reqR_unguarded(12) <= binary_1467_inst_req_1;
      reqR_unguarded(11) <= binary_1472_inst_req_1;
      reqR_unguarded(10) <= binary_1477_inst_req_1;
      reqR_unguarded(9) <= binary_1492_inst_req_1;
      reqR_unguarded(8) <= binary_1507_inst_req_1;
      reqR_unguarded(7) <= binary_1512_inst_req_1;
      reqR_unguarded(6) <= binary_1517_inst_req_1;
      reqR_unguarded(5) <= binary_1548_inst_req_1;
      reqR_unguarded(4) <= binary_1563_inst_req_1;
      reqR_unguarded(3) <= binary_1568_inst_req_1;
      reqR_unguarded(2) <= binary_1573_inst_req_1;
      reqR_unguarded(1) <= binary_1588_inst_req_1;
      reqR_unguarded(0) <= binary_1603_inst_req_1;
      binary_1844_inst_ack_1 <= ackR_unguarded(63);
      binary_1764_inst_ack_1 <= ackR_unguarded(62);
      binary_1608_inst_ack_1 <= ackR_unguarded(61);
      binary_1789_inst_ack_1 <= ackR_unguarded(60);
      binary_1784_inst_ack_1 <= ackR_unguarded(59);
      binary_1829_inst_ack_1 <= ackR_unguarded(58);
      binary_1859_inst_ack_1 <= ackR_unguarded(57);
      binary_1864_inst_ack_1 <= ackR_unguarded(56);
      binary_1824_inst_ack_1 <= ackR_unguarded(55);
      binary_1693_inst_ack_1 <= ackR_unguarded(54);
      binary_1819_inst_ack_1 <= ackR_unguarded(53);
      binary_1779_inst_ack_1 <= ackR_unguarded(52);
      binary_1869_inst_ack_1 <= ackR_unguarded(51);
      binary_1683_inst_ack_1 <= ackR_unguarded(50);
      binary_1628_inst_ack_1 <= ackR_unguarded(49);
      binary_1643_inst_ack_1 <= ackR_unguarded(48);
      binary_1613_inst_ack_1 <= ackR_unguarded(47);
      binary_1688_inst_ack_1 <= ackR_unguarded(46);
      binary_1648_inst_ack_1 <= ackR_unguarded(45);
      binary_1653_inst_ack_1 <= ackR_unguarded(44);
      binary_1724_inst_ack_1 <= ackR_unguarded(43);
      binary_1739_inst_ack_1 <= ackR_unguarded(42);
      binary_1744_inst_ack_1 <= ackR_unguarded(41);
      binary_1749_inst_ack_1 <= ackR_unguarded(40);
      binary_1668_inst_ack_1 <= ackR_unguarded(39);
      binary_1804_inst_ack_1 <= ackR_unguarded(38);
      binary_1148_inst_ack_1 <= ackR_unguarded(37);
      binary_1163_inst_ack_1 <= ackR_unguarded(36);
      binary_1168_inst_ack_1 <= ackR_unguarded(35);
      binary_1173_inst_ack_1 <= ackR_unguarded(34);
      binary_1204_inst_ack_1 <= ackR_unguarded(33);
      binary_1219_inst_ack_1 <= ackR_unguarded(32);
      binary_1224_inst_ack_1 <= ackR_unguarded(31);
      binary_1229_inst_ack_1 <= ackR_unguarded(30);
      binary_1260_inst_ack_1 <= ackR_unguarded(29);
      binary_1275_inst_ack_1 <= ackR_unguarded(28);
      binary_1280_inst_ack_1 <= ackR_unguarded(27);
      binary_1285_inst_ack_1 <= ackR_unguarded(26);
      binary_1316_inst_ack_1 <= ackR_unguarded(25);
      binary_1331_inst_ack_1 <= ackR_unguarded(24);
      binary_1336_inst_ack_1 <= ackR_unguarded(23);
      binary_1341_inst_ack_1 <= ackR_unguarded(22);
      binary_1372_inst_ack_1 <= ackR_unguarded(21);
      binary_1387_inst_ack_1 <= ackR_unguarded(20);
      binary_1392_inst_ack_1 <= ackR_unguarded(19);
      binary_1397_inst_ack_1 <= ackR_unguarded(18);
      binary_1412_inst_ack_1 <= ackR_unguarded(17);
      binary_1427_inst_ack_1 <= ackR_unguarded(16);
      binary_1432_inst_ack_1 <= ackR_unguarded(15);
      binary_1437_inst_ack_1 <= ackR_unguarded(14);
      binary_1452_inst_ack_1 <= ackR_unguarded(13);
      binary_1467_inst_ack_1 <= ackR_unguarded(12);
      binary_1472_inst_ack_1 <= ackR_unguarded(11);
      binary_1477_inst_ack_1 <= ackR_unguarded(10);
      binary_1492_inst_ack_1 <= ackR_unguarded(9);
      binary_1507_inst_ack_1 <= ackR_unguarded(8);
      binary_1512_inst_ack_1 <= ackR_unguarded(7);
      binary_1517_inst_ack_1 <= ackR_unguarded(6);
      binary_1548_inst_ack_1 <= ackR_unguarded(5);
      binary_1563_inst_ack_1 <= ackR_unguarded(4);
      binary_1568_inst_ack_1 <= ackR_unguarded(3);
      binary_1573_inst_ack_1 <= ackR_unguarded(2);
      binary_1588_inst_ack_1 <= ackR_unguarded(1);
      binary_1603_inst_ack_1 <= ackR_unguarded(0);
      gI0: GuardInterface generic map(nreqs => 64) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 64) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          operator_id => "ApFloatAdd",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 64 -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : binary_1875_inst 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_743;
      indvarx_xnext_1876 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_1875_inst_req_0;
      reqR(0) <= binary_1875_inst_req_1;
      binary_1875_inst_ack_0 <= ackL(0); 
      binary_1875_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : binary_1881_inst 
    ApIntEq_group_54: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xnext_1876;
      exitcond222_1882 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_1881_inst_req_0;
      reqR(0) <= binary_1881_inst_req_1;
      binary_1881_inst_ack_0 <= ackL(0); 
      binary_1881_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : binary_2023_inst 
    ApIntAdd_group_55: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar56_589;
      indvarx_xnext57_2024 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_2023_inst_req_0;
      reqR(0) <= binary_2023_inst_req_1;
      binary_2023_inst_ack_0 <= ackL(0); 
      binary_2023_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : binary_2029_inst 
    ApIntEq_group_56: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xnext57_2024;
      exitcond_2030 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_2029_inst_req_0;
      reqR(0) <= binary_2029_inst_req_1;
      binary_2029_inst_ack_0 <= ackL(0); 
      binary_2029_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : binary_2042_inst 
    ApIntAdd_group_57: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar60_555;
      indvarx_xnext61_2043 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_2042_inst_req_0;
      reqR(0) <= binary_2042_inst_req_1;
      binary_2042_inst_ack_0 <= ackL(0); 
      binary_2042_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : binary_2048_inst 
    ApIntEq_group_58: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xnext61_2043;
      exitcond310_2049 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_2048_inst_req_0;
      reqR(0) <= binary_2048_inst_req_1;
      binary_2048_inst_ack_0 <= ackL(0); 
      binary_2048_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : binary_987_inst binary_867_inst binary_567_inst binary_601_inst binary_721_inst 
    ApIntMul_group_59: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      -- 
    begin -- 
      data_in <= indvar_743 & indvar_743 & indvar60_555 & indvar56_589 & indvar56_589;
      tmp266_988 <= data_out(159 downto 128);
      tmp335_868 <= data_out(127 downto 96);
      tmp311_568 <= data_out(95 downto 64);
      tmp312_602 <= data_out(63 downto 32);
      tmp268_722 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      reqL_unguarded(4) <= binary_987_inst_req_0;
      reqL_unguarded(3) <= binary_867_inst_req_0;
      reqL_unguarded(2) <= binary_567_inst_req_0;
      reqL_unguarded(1) <= binary_601_inst_req_0;
      reqL_unguarded(0) <= binary_721_inst_req_0;
      binary_987_inst_ack_0 <= ackL_unguarded(4);
      binary_867_inst_ack_0 <= ackL_unguarded(3);
      binary_567_inst_ack_0 <= ackL_unguarded(2);
      binary_601_inst_ack_0 <= ackL_unguarded(1);
      binary_721_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= binary_987_inst_req_1;
      reqR_unguarded(3) <= binary_867_inst_req_1;
      reqR_unguarded(2) <= binary_567_inst_req_1;
      reqR_unguarded(1) <= binary_601_inst_req_1;
      reqR_unguarded(0) <= binary_721_inst_req_1;
      binary_987_inst_ack_1 <= ackR_unguarded(4);
      binary_867_inst_ack_1 <= ackR_unguarded(3);
      binary_567_inst_ack_1 <= ackR_unguarded(2);
      binary_601_inst_ack_1 <= ackR_unguarded(1);
      binary_721_inst_ack_1 <= ackR_unguarded(0);
      gI0: GuardInterface generic map(nreqs => 5) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 5) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 5--
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : binary_573_inst 
    ApIntAdd_group_60: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp311_568;
      tmp318_574 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_573_inst_req_0;
      reqR(0) <= binary_573_inst_req_1;
      binary_573_inst_ack_0 <= ackL(0); 
      binary_573_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : binary_579_inst 
    ApIntAdd_group_61: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp311_568;
      tmp324_580 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_579_inst_req_0;
      reqR(0) <= binary_579_inst_req_1;
      binary_579_inst_ack_0 <= ackL(0); 
      binary_579_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : binary_585_inst 
    ApIntAdd_group_62: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp311_568;
      tmp329_586 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_585_inst_req_0;
      reqR(0) <= binary_585_inst_req_1;
      binary_585_inst_ack_0 <= ackL(0); 
      binary_585_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : binary_613_inst 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp312_602;
      tmp314_614 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_613_inst_req_0;
      reqR(0) <= binary_613_inst_req_1;
      binary_613_inst_ack_0 <= ackL(0); 
      binary_613_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : binary_625_inst 
    ApIntAdd_group_64: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp312_602;
      tmp316_626 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_625_inst_req_0;
      reqR(0) <= binary_625_inst_req_1;
      binary_625_inst_ack_0 <= ackL(0); 
      binary_625_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : binary_655_inst 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp312_602;
      tmp322_656 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_655_inst_req_0;
      reqR(0) <= binary_655_inst_req_1;
      binary_655_inst_ack_0 <= ackL(0); 
      binary_655_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : binary_727_inst 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp268_722;
      tmp275_728 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_727_inst_req_0;
      reqR(0) <= binary_727_inst_req_1;
      binary_727_inst_ack_0 <= ackL(0); 
      binary_727_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : binary_733_inst 
    ApIntAdd_group_67: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp268_722;
      tmp280_734 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_733_inst_req_0;
      reqR(0) <= binary_733_inst_req_1;
      binary_733_inst_ack_0 <= ackL(0); 
      binary_733_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : binary_739_inst 
    ApIntAdd_group_68: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp268_722;
      tmp285_740 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_739_inst_req_0;
      reqR(0) <= binary_739_inst_req_1;
      binary_739_inst_ack_0 <= ackL(0); 
      binary_739_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : binary_879_inst 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp335_868;
      tmp337_880 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_879_inst_req_0;
      reqR(0) <= binary_879_inst_req_1;
      binary_879_inst_ack_0 <= ackL(0); 
      binary_879_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : binary_891_inst 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp335_868;
      tmp339_892 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_891_inst_req_0;
      reqR(0) <= binary_891_inst_req_1;
      binary_891_inst_ack_0 <= ackL(0); 
      binary_891_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : binary_921_inst 
    ApIntAdd_group_71: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp335_868;
      tmp344_922 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_921_inst_req_0;
      reqR(0) <= binary_921_inst_req_1;
      binary_921_inst_ack_0 <= ackL(0); 
      binary_921_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : binary_993_inst 
    ApIntAdd_group_72: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp266_988;
      tmp267_994 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_993_inst_req_0;
      reqR(0) <= binary_993_inst_req_1;
      binary_993_inst_ack_0 <= ackL(0); 
      binary_993_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared load operator group (0) : ptr_deref_1697_load_0 ptr_deref_1701_load_0 ptr_deref_1709_load_0 ptr_deref_1705_load_0 ptr_deref_1105_load_0 ptr_deref_1113_load_0 ptr_deref_1121_load_0 ptr_deref_1129_load_0 ptr_deref_1345_load_0 ptr_deref_1349_load_0 ptr_deref_1353_load_0 ptr_deref_1357_load_0 ptr_deref_1521_load_0 ptr_deref_1525_load_0 ptr_deref_1529_load_0 ptr_deref_1533_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(143 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_1697_load_0_req_0;
      reqL_unguarded(14) <= ptr_deref_1701_load_0_req_0;
      reqL_unguarded(13) <= ptr_deref_1709_load_0_req_0;
      reqL_unguarded(12) <= ptr_deref_1705_load_0_req_0;
      reqL_unguarded(11) <= ptr_deref_1105_load_0_req_0;
      reqL_unguarded(10) <= ptr_deref_1113_load_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1121_load_0_req_0;
      reqL_unguarded(8) <= ptr_deref_1129_load_0_req_0;
      reqL_unguarded(7) <= ptr_deref_1345_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_1349_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_1353_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1357_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_1521_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1525_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1529_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1533_load_0_req_0;
      ptr_deref_1697_load_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_1701_load_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_1709_load_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_1705_load_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_1105_load_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_1113_load_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1121_load_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_1129_load_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_1345_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_1349_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_1353_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1357_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_1521_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1525_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1529_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1533_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_1697_load_0_req_1;
      reqR_unguarded(14) <= ptr_deref_1701_load_0_req_1;
      reqR_unguarded(13) <= ptr_deref_1709_load_0_req_1;
      reqR_unguarded(12) <= ptr_deref_1705_load_0_req_1;
      reqR_unguarded(11) <= ptr_deref_1105_load_0_req_1;
      reqR_unguarded(10) <= ptr_deref_1113_load_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1121_load_0_req_1;
      reqR_unguarded(8) <= ptr_deref_1129_load_0_req_1;
      reqR_unguarded(7) <= ptr_deref_1345_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_1349_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_1353_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1357_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_1521_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1525_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1529_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1533_load_0_req_1;
      ptr_deref_1697_load_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_1701_load_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_1709_load_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_1705_load_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_1105_load_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_1113_load_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1121_load_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_1129_load_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_1345_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_1349_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_1353_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1357_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_1521_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1525_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1529_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1533_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 16) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 16) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1697_word_address_0 & ptr_deref_1701_word_address_0 & ptr_deref_1709_word_address_0 & ptr_deref_1705_word_address_0 & ptr_deref_1105_word_address_0 & ptr_deref_1113_word_address_0 & ptr_deref_1121_word_address_0 & ptr_deref_1129_word_address_0 & ptr_deref_1345_word_address_0 & ptr_deref_1349_word_address_0 & ptr_deref_1353_word_address_0 & ptr_deref_1357_word_address_0 & ptr_deref_1521_word_address_0 & ptr_deref_1525_word_address_0 & ptr_deref_1529_word_address_0 & ptr_deref_1533_word_address_0;
      ptr_deref_1697_data_0 <= data_out(511 downto 480);
      ptr_deref_1701_data_0 <= data_out(479 downto 448);
      ptr_deref_1709_data_0 <= data_out(447 downto 416);
      ptr_deref_1705_data_0 <= data_out(415 downto 384);
      ptr_deref_1105_data_0 <= data_out(383 downto 352);
      ptr_deref_1113_data_0 <= data_out(351 downto 320);
      ptr_deref_1121_data_0 <= data_out(319 downto 288);
      ptr_deref_1129_data_0 <= data_out(287 downto 256);
      ptr_deref_1345_data_0 <= data_out(255 downto 224);
      ptr_deref_1349_data_0 <= data_out(223 downto 192);
      ptr_deref_1353_data_0 <= data_out(191 downto 160);
      ptr_deref_1357_data_0 <= data_out(159 downto 128);
      ptr_deref_1521_data_0 <= data_out(127 downto 96);
      ptr_deref_1525_data_0 <= data_out(95 downto 64);
      ptr_deref_1529_data_0 <= data_out(63 downto 32);
      ptr_deref_1533_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 9,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(8 downto 0),
          mtag => memory_space_0_lr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 16,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1109_load_0 ptr_deref_1117_load_0 ptr_deref_1125_load_0 ptr_deref_1133_load_0 ptr_deref_1177_load_0 ptr_deref_1181_load_0 ptr_deref_1185_load_0 ptr_deref_1189_load_0 ptr_deref_1233_load_0 ptr_deref_1237_load_0 ptr_deref_1241_load_0 ptr_deref_1245_load_0 ptr_deref_1289_load_0 ptr_deref_1293_load_0 ptr_deref_1297_load_0 ptr_deref_1301_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(143 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_1109_load_0_req_0;
      reqL_unguarded(14) <= ptr_deref_1117_load_0_req_0;
      reqL_unguarded(13) <= ptr_deref_1125_load_0_req_0;
      reqL_unguarded(12) <= ptr_deref_1133_load_0_req_0;
      reqL_unguarded(11) <= ptr_deref_1177_load_0_req_0;
      reqL_unguarded(10) <= ptr_deref_1181_load_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1185_load_0_req_0;
      reqL_unguarded(8) <= ptr_deref_1189_load_0_req_0;
      reqL_unguarded(7) <= ptr_deref_1233_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_1237_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_1241_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1245_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_1289_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1293_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1297_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1301_load_0_req_0;
      ptr_deref_1109_load_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_1117_load_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_1125_load_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_1133_load_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_1177_load_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_1181_load_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1185_load_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_1189_load_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_1233_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_1237_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_1241_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1245_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_1289_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1293_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1297_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1301_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_1109_load_0_req_1;
      reqR_unguarded(14) <= ptr_deref_1117_load_0_req_1;
      reqR_unguarded(13) <= ptr_deref_1125_load_0_req_1;
      reqR_unguarded(12) <= ptr_deref_1133_load_0_req_1;
      reqR_unguarded(11) <= ptr_deref_1177_load_0_req_1;
      reqR_unguarded(10) <= ptr_deref_1181_load_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1185_load_0_req_1;
      reqR_unguarded(8) <= ptr_deref_1189_load_0_req_1;
      reqR_unguarded(7) <= ptr_deref_1233_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_1237_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_1241_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1245_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_1289_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1293_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1297_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1301_load_0_req_1;
      ptr_deref_1109_load_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_1117_load_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_1125_load_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_1133_load_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_1177_load_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_1181_load_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1185_load_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_1189_load_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_1233_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_1237_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_1241_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1245_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_1289_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1293_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1297_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1301_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 16) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 16) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1109_word_address_0 & ptr_deref_1117_word_address_0 & ptr_deref_1125_word_address_0 & ptr_deref_1133_word_address_0 & ptr_deref_1177_word_address_0 & ptr_deref_1181_word_address_0 & ptr_deref_1185_word_address_0 & ptr_deref_1189_word_address_0 & ptr_deref_1233_word_address_0 & ptr_deref_1237_word_address_0 & ptr_deref_1241_word_address_0 & ptr_deref_1245_word_address_0 & ptr_deref_1289_word_address_0 & ptr_deref_1293_word_address_0 & ptr_deref_1297_word_address_0 & ptr_deref_1301_word_address_0;
      ptr_deref_1109_data_0 <= data_out(511 downto 480);
      ptr_deref_1117_data_0 <= data_out(479 downto 448);
      ptr_deref_1125_data_0 <= data_out(447 downto 416);
      ptr_deref_1133_data_0 <= data_out(415 downto 384);
      ptr_deref_1177_data_0 <= data_out(383 downto 352);
      ptr_deref_1181_data_0 <= data_out(351 downto 320);
      ptr_deref_1185_data_0 <= data_out(319 downto 288);
      ptr_deref_1189_data_0 <= data_out(287 downto 256);
      ptr_deref_1233_data_0 <= data_out(255 downto 224);
      ptr_deref_1237_data_0 <= data_out(223 downto 192);
      ptr_deref_1241_data_0 <= data_out(191 downto 160);
      ptr_deref_1245_data_0 <= data_out(159 downto 128);
      ptr_deref_1289_data_0 <= data_out(127 downto 96);
      ptr_deref_1293_data_0 <= data_out(95 downto 64);
      ptr_deref_1297_data_0 <= data_out(63 downto 32);
      ptr_deref_1301_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 9,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(8 downto 0),
          mtag => memory_space_1_lr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 16,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_1968_store_0 ptr_deref_2000_store_0 ptr_deref_2008_store_0 ptr_deref_2016_store_0 ptr_deref_1964_store_0 ptr_deref_2012_store_0 ptr_deref_1972_store_0 ptr_deref_1976_store_0 ptr_deref_1980_store_0 ptr_deref_1984_store_0 ptr_deref_1988_store_0 ptr_deref_1992_store_0 ptr_deref_1956_store_0 ptr_deref_2004_store_0 ptr_deref_1996_store_0 ptr_deref_1960_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(143 downto 0);
      signal data_in: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_1968_store_0_req_0;
      reqL_unguarded(14) <= ptr_deref_2000_store_0_req_0;
      reqL_unguarded(13) <= ptr_deref_2008_store_0_req_0;
      reqL_unguarded(12) <= ptr_deref_2016_store_0_req_0;
      reqL_unguarded(11) <= ptr_deref_1964_store_0_req_0;
      reqL_unguarded(10) <= ptr_deref_2012_store_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1972_store_0_req_0;
      reqL_unguarded(8) <= ptr_deref_1976_store_0_req_0;
      reqL_unguarded(7) <= ptr_deref_1980_store_0_req_0;
      reqL_unguarded(6) <= ptr_deref_1984_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_1988_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1992_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_1956_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_2004_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1996_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1960_store_0_req_0;
      ptr_deref_1968_store_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_2000_store_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_2008_store_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_2016_store_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_1964_store_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_2012_store_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1972_store_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_1976_store_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_1980_store_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_1984_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_1988_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1992_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_1956_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_2004_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1996_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1960_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_1968_store_0_req_1;
      reqR_unguarded(14) <= ptr_deref_2000_store_0_req_1;
      reqR_unguarded(13) <= ptr_deref_2008_store_0_req_1;
      reqR_unguarded(12) <= ptr_deref_2016_store_0_req_1;
      reqR_unguarded(11) <= ptr_deref_1964_store_0_req_1;
      reqR_unguarded(10) <= ptr_deref_2012_store_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1972_store_0_req_1;
      reqR_unguarded(8) <= ptr_deref_1976_store_0_req_1;
      reqR_unguarded(7) <= ptr_deref_1980_store_0_req_1;
      reqR_unguarded(6) <= ptr_deref_1984_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_1988_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1992_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_1956_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_2004_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1996_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1960_store_0_req_1;
      ptr_deref_1968_store_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_2000_store_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_2008_store_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_2016_store_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_1964_store_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_2012_store_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1972_store_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_1976_store_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_1980_store_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_1984_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_1988_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1992_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_1956_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_2004_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1996_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1960_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 16) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL,
        ackR => ackL,
        guards => guard_vector); -- 
      gI1: GuardInterface generic map(nreqs => 16) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1968_word_address_0 & ptr_deref_2000_word_address_0 & ptr_deref_2008_word_address_0 & ptr_deref_2016_word_address_0 & ptr_deref_1964_word_address_0 & ptr_deref_2012_word_address_0 & ptr_deref_1972_word_address_0 & ptr_deref_1976_word_address_0 & ptr_deref_1980_word_address_0 & ptr_deref_1984_word_address_0 & ptr_deref_1988_word_address_0 & ptr_deref_1992_word_address_0 & ptr_deref_1956_word_address_0 & ptr_deref_2004_word_address_0 & ptr_deref_1996_word_address_0 & ptr_deref_1960_word_address_0;
      data_in <= ptr_deref_1968_data_0 & ptr_deref_2000_data_0 & ptr_deref_2008_data_0 & ptr_deref_2016_data_0 & ptr_deref_1964_data_0 & ptr_deref_2012_data_0 & ptr_deref_1972_data_0 & ptr_deref_1976_data_0 & ptr_deref_1980_data_0 & ptr_deref_1984_data_0 & ptr_deref_1988_data_0 & ptr_deref_1992_data_0 & ptr_deref_1956_data_0 & ptr_deref_2004_data_0 & ptr_deref_1996_data_0 & ptr_deref_1960_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 9,
        data_width => 32,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(8 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 16,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    result_pipe_pipe_read_data: out std_logic_vector(31 downto 0);
    result_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    result_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(8 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(7 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(7 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(8 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(7 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module mmultiply
  component mmultiply is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
      in_data_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      result_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      result_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      result_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      mmultiply_base_call_reqs : out  std_logic_vector(0 downto 0);
      mmultiply_base_call_acks : in   std_logic_vector(0 downto 0);
      mmultiply_base_call_tag  :  out  std_logic_vector(0 downto 0);
      mmultiply_base_return_reqs : out  std_logic_vector(0 downto 0);
      mmultiply_base_return_acks : in   std_logic_vector(0 downto 0);
      mmultiply_base_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module mmultiply
  signal mmultiply_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal mmultiply_tag_out   : std_logic_vector(1 downto 0);
  signal mmultiply_start_req : std_logic;
  signal mmultiply_start_ack : std_logic;
  signal mmultiply_fin_req   : std_logic;
  signal mmultiply_fin_ack : std_logic;
  -- declarations related to module mmultiply_base
  component mmultiply_base is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module mmultiply_base
  signal mmultiply_base_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal mmultiply_base_tag_out   : std_logic_vector(1 downto 0);
  signal mmultiply_base_start_req : std_logic;
  signal mmultiply_base_start_ack : std_logic;
  signal mmultiply_base_fin_req   : std_logic;
  signal mmultiply_base_fin_ack : std_logic;
  -- caller side aggregated signals for module mmultiply_base
  signal mmultiply_base_call_reqs: std_logic_vector(0 downto 0);
  signal mmultiply_base_call_acks: std_logic_vector(0 downto 0);
  signal mmultiply_base_return_reqs: std_logic_vector(0 downto 0);
  signal mmultiply_base_return_acks: std_logic_vector(0 downto 0);
  signal mmultiply_base_call_tag: std_logic_vector(0 downto 0);
  signal mmultiply_base_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_pipe
  signal in_data_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe result_pipe
  signal result_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal result_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal result_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module mmultiply
  mmultiply_instance:mmultiply-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => mmultiply_start_req,
      start_ack => mmultiply_start_ack,
      fin_req => mmultiply_fin_req,
      fin_ack => mmultiply_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(8 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(7 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(4 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(8 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(7 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(4 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(8 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(7 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(4 downto 0),
      in_data_pipe_pipe_read_req => in_data_pipe_pipe_read_req(0 downto 0),
      in_data_pipe_pipe_read_ack => in_data_pipe_pipe_read_ack(0 downto 0),
      in_data_pipe_pipe_read_data => in_data_pipe_pipe_read_data(31 downto 0),
      result_pipe_pipe_write_req => result_pipe_pipe_write_req(0 downto 0),
      result_pipe_pipe_write_ack => result_pipe_pipe_write_ack(0 downto 0),
      result_pipe_pipe_write_data => result_pipe_pipe_write_data(31 downto 0),
      mmultiply_base_call_reqs => mmultiply_base_call_reqs(0 downto 0),
      mmultiply_base_call_acks => mmultiply_base_call_acks(0 downto 0),
      mmultiply_base_call_tag => mmultiply_base_call_tag(0 downto 0),
      mmultiply_base_return_reqs => mmultiply_base_return_reqs(0 downto 0),
      mmultiply_base_return_acks => mmultiply_base_return_acks(0 downto 0),
      mmultiply_base_return_tag => mmultiply_base_return_tag(0 downto 0),
      tag_in => mmultiply_tag_in,
      tag_out => mmultiply_tag_out-- 
    ); -- 
  -- module will be run forever 
  mmultiply_tag_in <= (others => '0');
  mmultiply_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => mmultiply_start_req, start_ack => mmultiply_start_ack,  fin_req => mmultiply_fin_req,  fin_ack => mmultiply_fin_ack);
  -- module mmultiply_base
  -- call arbiter for module mmultiply_base
  mmultiply_base_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => mmultiply_base_call_reqs,
      call_acks => mmultiply_base_call_acks,
      return_reqs => mmultiply_base_return_reqs,
      return_acks => mmultiply_base_return_acks,
      call_tag  => mmultiply_base_call_tag,
      return_tag  => mmultiply_base_return_tag,
      call_mtag => mmultiply_base_tag_in,
      return_mtag => mmultiply_base_tag_out,
      call_mreq => mmultiply_base_start_req,
      call_mack => mmultiply_base_start_ack,
      return_mreq => mmultiply_base_fin_req,
      return_mack => mmultiply_base_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  mmultiply_base_instance:mmultiply_base-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => mmultiply_base_start_req,
      start_ack => mmultiply_base_start_ack,
      fin_req => mmultiply_base_fin_req,
      fin_ack => mmultiply_base_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(8 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(7 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(4 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(8 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(7 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(4 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(8 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(7 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 0),
      tag_in => mmultiply_base_tag_in,
      tag_out => mmultiply_base_tag_out-- 
    ); -- 
  in_data_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_pipe_read_req,
      read_ack => in_data_pipe_pipe_read_ack,
      read_data => in_data_pipe_pipe_read_data,
      write_req => in_data_pipe_pipe_write_req,
      write_ack => in_data_pipe_pipe_write_ack,
      write_data => in_data_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  result_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => result_pipe_pipe_read_req,
      read_ack => result_pipe_pipe_read_ack,
      read_data => result_pipe_pipe_read_data,
      write_req => result_pipe_pipe_write_req,
      write_ack => result_pipe_pipe_write_ack,
      write_data => result_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 9,
      data_width => 32,
      tag_width => 5,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 9,
      data_width => 32,
      tag_width => 5,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 9,
      data_width => 32,
      tag_width => 5,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
