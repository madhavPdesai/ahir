-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant free_list_base_address : std_logic_vector(2 downto 0) := "000";
  constant head_base_address : std_logic_vector(0 downto 0) := "0";
  constant mempool_base_address : std_logic_vector(0 downto 0) := "0";
  constant xx_xstr1_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr2_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr3_base_address : std_logic_vector(2 downto 0) := "000";
  constant xx_xstr4_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr5_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr6_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr_base_address : std_logic_vector(4 downto 0) := "00000";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity foo is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    foo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
    foo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
    foo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
    foo_out_pipe_write_req : out  std_logic_vector(0 downto 0);
    foo_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
    foo_out_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity foo;
architecture Default of foo is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_89_root_address_inst_req_0 : boolean;
  signal array_obj_ref_89_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_89_root_address_inst_req_1 : boolean;
  signal array_obj_ref_89_root_address_inst_ack_1 : boolean;
  signal simple_obj_ref_71_inst_req_0 : boolean;
  signal simple_obj_ref_71_inst_ack_0 : boolean;
  signal type_cast_72_inst_req_0 : boolean;
  signal type_cast_72_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal ptr_deref_79_gather_scatter_req_0 : boolean;
  signal ptr_deref_79_gather_scatter_ack_0 : boolean;
  signal ptr_deref_79_store_0_req_0 : boolean;
  signal ptr_deref_79_store_0_ack_0 : boolean;
  signal ptr_deref_79_store_0_req_1 : boolean;
  signal ptr_deref_79_store_0_ack_1 : boolean;
  signal ptr_deref_84_load_0_req_0 : boolean;
  signal ptr_deref_84_load_0_ack_0 : boolean;
  signal ptr_deref_84_load_0_req_1 : boolean;
  signal ptr_deref_84_load_0_ack_1 : boolean;
  signal ptr_deref_84_gather_scatter_req_0 : boolean;
  signal ptr_deref_84_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_89_base_resize_req_0 : boolean;
  signal array_obj_ref_89_base_resize_ack_0 : boolean;
  signal type_cast_119_inst_req_0 : boolean;
  signal type_cast_119_inst_ack_0 : boolean;
  signal array_obj_ref_89_final_reg_req_0 : boolean;
  signal array_obj_ref_89_final_reg_ack_0 : boolean;
  signal ptr_deref_93_base_resize_req_0 : boolean;
  signal ptr_deref_93_base_resize_ack_0 : boolean;
  signal ptr_deref_93_root_address_inst_req_0 : boolean;
  signal ptr_deref_93_root_address_inst_ack_0 : boolean;
  signal ptr_deref_93_addr_0_req_0 : boolean;
  signal ptr_deref_93_addr_0_ack_0 : boolean;
  signal ptr_deref_93_load_0_req_0 : boolean;
  signal ptr_deref_93_load_0_ack_0 : boolean;
  signal ptr_deref_93_load_0_req_1 : boolean;
  signal ptr_deref_93_load_0_ack_1 : boolean;
  signal ptr_deref_93_gather_scatter_req_0 : boolean;
  signal ptr_deref_93_gather_scatter_ack_0 : boolean;
  signal binary_98_inst_req_0 : boolean;
  signal binary_98_inst_ack_0 : boolean;
  signal binary_98_inst_req_1 : boolean;
  signal binary_98_inst_ack_1 : boolean;
  signal ptr_deref_102_load_0_req_0 : boolean;
  signal ptr_deref_102_load_0_ack_0 : boolean;
  signal ptr_deref_102_load_0_req_1 : boolean;
  signal ptr_deref_102_load_0_ack_1 : boolean;
  signal ptr_deref_102_gather_scatter_req_0 : boolean;
  signal ptr_deref_102_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_107_base_resize_req_0 : boolean;
  signal array_obj_ref_107_base_resize_ack_0 : boolean;
  signal array_obj_ref_107_root_address_inst_req_0 : boolean;
  signal array_obj_ref_107_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_107_root_address_inst_req_1 : boolean;
  signal array_obj_ref_107_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_107_final_reg_req_0 : boolean;
  signal array_obj_ref_107_final_reg_ack_0 : boolean;
  signal ptr_deref_110_base_resize_req_0 : boolean;
  signal ptr_deref_110_base_resize_ack_0 : boolean;
  signal ptr_deref_110_root_address_inst_req_0 : boolean;
  signal ptr_deref_110_root_address_inst_ack_0 : boolean;
  signal ptr_deref_110_addr_0_req_0 : boolean;
  signal ptr_deref_110_addr_0_ack_0 : boolean;
  signal ptr_deref_110_gather_scatter_req_0 : boolean;
  signal ptr_deref_110_gather_scatter_ack_0 : boolean;
  signal ptr_deref_110_store_0_req_0 : boolean;
  signal ptr_deref_110_store_0_ack_0 : boolean;
  signal ptr_deref_110_store_0_req_1 : boolean;
  signal ptr_deref_110_store_0_ack_1 : boolean;
  signal ptr_deref_115_load_0_req_0 : boolean;
  signal ptr_deref_115_load_0_ack_0 : boolean;
  signal ptr_deref_115_load_0_req_1 : boolean;
  signal ptr_deref_115_load_0_ack_1 : boolean;
  signal ptr_deref_115_gather_scatter_req_0 : boolean;
  signal ptr_deref_115_gather_scatter_ack_0 : boolean;
  signal type_cast_128_inst_req_0 : boolean;
  signal type_cast_128_inst_ack_0 : boolean;
  signal simple_obj_ref_126_inst_req_0 : boolean;
  signal simple_obj_ref_126_inst_ack_0 : boolean;
  signal memory_space_10_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_10_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_10_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_10_lr_tag : std_logic_vector(2 downto 0);
  signal memory_space_10_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_10_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_10_lc_data : std_logic_vector(95 downto 0);
  signal memory_space_10_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_10_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_10_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  foo_CP_0: Block -- control-path 
    signal foo_CP_0_start: Boolean;
    signal Xentry_1_symbol: Boolean;
    signal Xexit_2_symbol: Boolean;
    signal branch_block_stmt_56_3_symbol : Boolean;
    -- 
  begin -- 
    foo_CP_0_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_1_symbol  <= foo_CP_0_start; -- transition $entry
    branch_block_stmt_56_3: Block -- branch_block_stmt_56 
      signal branch_block_stmt_56_3_start: Boolean;
      signal Xentry_4_symbol: Boolean;
      signal Xexit_5_symbol: Boolean;
      signal branch_block_stmt_56_x_xentry_x_xx_x6_symbol : Boolean;
      signal branch_block_stmt_56_x_xexit_x_xx_x7_symbol : Boolean;
      signal assign_stmt_61_x_xentry_x_xx_x8_symbol : Boolean;
      signal assign_stmt_61_x_xexit_x_xx_x9_symbol : Boolean;
      signal bb_0_bb_1_10_symbol : Boolean;
      signal merge_stmt_63_x_xexit_x_xx_x11_symbol : Boolean;
      signal assign_stmt_68_x_xentry_x_xx_x12_symbol : Boolean;
      signal assign_stmt_68_x_xexit_x_xx_x13_symbol : Boolean;
      signal assign_stmt_73_x_xentry_x_xx_x14_symbol : Boolean;
      signal assign_stmt_73_x_xexit_x_xx_x15_symbol : Boolean;
      signal assign_stmt_77_to_assign_stmt_125_x_xentry_x_xx_x16_symbol : Boolean;
      signal assign_stmt_77_to_assign_stmt_125_x_xexit_x_xx_x17_symbol : Boolean;
      signal assign_stmt_129_x_xentry_x_xx_x18_symbol : Boolean;
      signal assign_stmt_129_x_xexit_x_xx_x19_symbol : Boolean;
      signal bb_1_bb_1_20_symbol : Boolean;
      signal assign_stmt_61_21_symbol : Boolean;
      signal assign_stmt_68_24_symbol : Boolean;
      signal assign_stmt_73_27_symbol : Boolean;
      signal assign_stmt_77_to_assign_stmt_125_45_symbol : Boolean;
      signal assign_stmt_129_352_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_371_symbol : Boolean;
      signal bb_1_bb_1_PhiReq_374_symbol : Boolean;
      signal merge_stmt_63_PhiReqMerge_377_symbol : Boolean;
      signal merge_stmt_63_PhiAck_378_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_56_3_start <= Xentry_1_symbol; -- control passed to block
      Xentry_4_symbol  <= branch_block_stmt_56_3_start; -- transition branch_block_stmt_56/$entry
      branch_block_stmt_56_x_xentry_x_xx_x6_symbol  <=  Xentry_4_symbol; -- place branch_block_stmt_56/branch_block_stmt_56__entry__ (optimized away) 
      branch_block_stmt_56_x_xexit_x_xx_x7_symbol  <=   false ; -- place branch_block_stmt_56/branch_block_stmt_56__exit__ (optimized away) 
      assign_stmt_61_x_xentry_x_xx_x8_symbol  <=  branch_block_stmt_56_x_xentry_x_xx_x6_symbol; -- place branch_block_stmt_56/assign_stmt_61__entry__ (optimized away) 
      assign_stmt_61_x_xexit_x_xx_x9_symbol  <=  assign_stmt_61_21_symbol; -- place branch_block_stmt_56/assign_stmt_61__exit__ (optimized away) 
      bb_0_bb_1_10_symbol  <=  assign_stmt_61_x_xexit_x_xx_x9_symbol; -- place branch_block_stmt_56/bb_0_bb_1 (optimized away) 
      merge_stmt_63_x_xexit_x_xx_x11_symbol  <=  merge_stmt_63_PhiAck_378_symbol; -- place branch_block_stmt_56/merge_stmt_63__exit__ (optimized away) 
      assign_stmt_68_x_xentry_x_xx_x12_symbol  <=  merge_stmt_63_x_xexit_x_xx_x11_symbol; -- place branch_block_stmt_56/assign_stmt_68__entry__ (optimized away) 
      assign_stmt_68_x_xexit_x_xx_x13_symbol  <=  assign_stmt_68_24_symbol; -- place branch_block_stmt_56/assign_stmt_68__exit__ (optimized away) 
      assign_stmt_73_x_xentry_x_xx_x14_symbol  <=  assign_stmt_68_x_xexit_x_xx_x13_symbol; -- place branch_block_stmt_56/assign_stmt_73__entry__ (optimized away) 
      assign_stmt_73_x_xexit_x_xx_x15_symbol  <=  assign_stmt_73_27_symbol; -- place branch_block_stmt_56/assign_stmt_73__exit__ (optimized away) 
      assign_stmt_77_to_assign_stmt_125_x_xentry_x_xx_x16_symbol  <=  assign_stmt_73_x_xexit_x_xx_x15_symbol; -- place branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125__entry__ (optimized away) 
      assign_stmt_77_to_assign_stmt_125_x_xexit_x_xx_x17_symbol  <=  assign_stmt_77_to_assign_stmt_125_45_symbol; -- place branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125__exit__ (optimized away) 
      assign_stmt_129_x_xentry_x_xx_x18_symbol  <=  assign_stmt_77_to_assign_stmt_125_x_xexit_x_xx_x17_symbol; -- place branch_block_stmt_56/assign_stmt_129__entry__ (optimized away) 
      assign_stmt_129_x_xexit_x_xx_x19_symbol  <=  assign_stmt_129_352_symbol; -- place branch_block_stmt_56/assign_stmt_129__exit__ (optimized away) 
      bb_1_bb_1_20_symbol  <=  assign_stmt_129_x_xexit_x_xx_x19_symbol; -- place branch_block_stmt_56/bb_1_bb_1 (optimized away) 
      assign_stmt_61_21: Block -- branch_block_stmt_56/assign_stmt_61 
        signal assign_stmt_61_21_start: Boolean;
        signal Xentry_22_symbol: Boolean;
        signal Xexit_23_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_61_21_start <= assign_stmt_61_x_xentry_x_xx_x8_symbol; -- control passed to block
        Xentry_22_symbol  <= assign_stmt_61_21_start; -- transition branch_block_stmt_56/assign_stmt_61/$entry
        Xexit_23_symbol <= Xentry_22_symbol; -- transition branch_block_stmt_56/assign_stmt_61/$exit
        assign_stmt_61_21_symbol <= Xexit_23_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_61
      assign_stmt_68_24: Block -- branch_block_stmt_56/assign_stmt_68 
        signal assign_stmt_68_24_start: Boolean;
        signal Xentry_25_symbol: Boolean;
        signal Xexit_26_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_68_24_start <= assign_stmt_68_x_xentry_x_xx_x12_symbol; -- control passed to block
        Xentry_25_symbol  <= assign_stmt_68_24_start; -- transition branch_block_stmt_56/assign_stmt_68/$entry
        Xexit_26_symbol <= Xentry_25_symbol; -- transition branch_block_stmt_56/assign_stmt_68/$exit
        assign_stmt_68_24_symbol <= Xexit_26_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_68
      assign_stmt_73_27: Block -- branch_block_stmt_56/assign_stmt_73 
        signal assign_stmt_73_27_start: Boolean;
        signal Xentry_28_symbol: Boolean;
        signal Xexit_29_symbol: Boolean;
        signal assign_stmt_73_active_x_x30_symbol : Boolean;
        signal assign_stmt_73_completed_x_x31_symbol : Boolean;
        signal type_cast_72_active_x_x32_symbol : Boolean;
        signal type_cast_72_trigger_x_x33_symbol : Boolean;
        signal simple_obj_ref_71_trigger_x_x34_symbol : Boolean;
        signal simple_obj_ref_71_complete_35_symbol : Boolean;
        signal type_cast_72_complete_40_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_73_27_start <= assign_stmt_73_x_xentry_x_xx_x14_symbol; -- control passed to block
        Xentry_28_symbol  <= assign_stmt_73_27_start; -- transition branch_block_stmt_56/assign_stmt_73/$entry
        assign_stmt_73_active_x_x30_symbol <= type_cast_72_complete_40_symbol; -- transition branch_block_stmt_56/assign_stmt_73/assign_stmt_73_active_
        assign_stmt_73_completed_x_x31_symbol <= assign_stmt_73_active_x_x30_symbol; -- transition branch_block_stmt_56/assign_stmt_73/assign_stmt_73_completed_
        type_cast_72_active_x_x32_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_73/type_cast_72_active_ 
          signal type_cast_72_active_x_x32_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_72_active_x_x32_predecessors(0) <= type_cast_72_trigger_x_x33_symbol;
          type_cast_72_active_x_x32_predecessors(1) <= simple_obj_ref_71_complete_35_symbol;
          type_cast_72_active_x_x32_join: join -- 
            port map( -- 
              preds => type_cast_72_active_x_x32_predecessors,
              symbol_out => type_cast_72_active_x_x32_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_73/type_cast_72_active_
        type_cast_72_trigger_x_x33_symbol <= Xentry_28_symbol; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_trigger_
        simple_obj_ref_71_trigger_x_x34_symbol <= Xentry_28_symbol; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_trigger_
        simple_obj_ref_71_complete_35: Block -- branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete 
          signal simple_obj_ref_71_complete_35_start: Boolean;
          signal Xentry_36_symbol: Boolean;
          signal Xexit_37_symbol: Boolean;
          signal req_38_symbol : Boolean;
          signal ack_39_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_71_complete_35_start <= simple_obj_ref_71_trigger_x_x34_symbol; -- control passed to block
          Xentry_36_symbol  <= simple_obj_ref_71_complete_35_start; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/$entry
          req_38_symbol <= Xentry_36_symbol; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/req
          simple_obj_ref_71_inst_req_0 <= req_38_symbol; -- link to DP
          ack_39_symbol <= simple_obj_ref_71_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/ack
          Xexit_37_symbol <= ack_39_symbol; -- transition branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete/$exit
          simple_obj_ref_71_complete_35_symbol <= Xexit_37_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_73/simple_obj_ref_71_complete
        type_cast_72_complete_40: Block -- branch_block_stmt_56/assign_stmt_73/type_cast_72_complete 
          signal type_cast_72_complete_40_start: Boolean;
          signal Xentry_41_symbol: Boolean;
          signal Xexit_42_symbol: Boolean;
          signal req_43_symbol : Boolean;
          signal ack_44_symbol : Boolean;
          -- 
        begin -- 
          type_cast_72_complete_40_start <= type_cast_72_active_x_x32_symbol; -- control passed to block
          Xentry_41_symbol  <= type_cast_72_complete_40_start; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/$entry
          req_43_symbol <= Xentry_41_symbol; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/req
          type_cast_72_inst_req_0 <= req_43_symbol; -- link to DP
          ack_44_symbol <= type_cast_72_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/ack
          Xexit_42_symbol <= ack_44_symbol; -- transition branch_block_stmt_56/assign_stmt_73/type_cast_72_complete/$exit
          type_cast_72_complete_40_symbol <= Xexit_42_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_73/type_cast_72_complete
        Xexit_29_symbol <= assign_stmt_73_completed_x_x31_symbol; -- transition branch_block_stmt_56/assign_stmt_73/$exit
        assign_stmt_73_27_symbol <= Xexit_29_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_73
      assign_stmt_77_to_assign_stmt_125_45: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125 
        signal assign_stmt_77_to_assign_stmt_125_45_start: Boolean;
        signal Xentry_46_symbol: Boolean;
        signal Xexit_47_symbol: Boolean;
        signal assign_stmt_77_active_x_x48_symbol : Boolean;
        signal assign_stmt_77_completed_x_x49_symbol : Boolean;
        signal type_cast_76_active_x_x50_symbol : Boolean;
        signal type_cast_76_trigger_x_x51_symbol : Boolean;
        signal simple_obj_ref_75_complete_52_symbol : Boolean;
        signal type_cast_76_complete_53_symbol : Boolean;
        signal assign_stmt_81_active_x_x58_symbol : Boolean;
        signal assign_stmt_81_completed_x_x59_symbol : Boolean;
        signal simple_obj_ref_80_complete_60_symbol : Boolean;
        signal ptr_deref_79_trigger_x_x61_symbol : Boolean;
        signal ptr_deref_79_active_x_x62_symbol : Boolean;
        signal ptr_deref_79_base_address_calculated_63_symbol : Boolean;
        signal ptr_deref_79_root_address_calculated_64_symbol : Boolean;
        signal ptr_deref_79_word_address_calculated_65_symbol : Boolean;
        signal ptr_deref_79_request_66_symbol : Boolean;
        signal ptr_deref_79_complete_79_symbol : Boolean;
        signal assign_stmt_85_active_x_x90_symbol : Boolean;
        signal assign_stmt_85_completed_x_x91_symbol : Boolean;
        signal ptr_deref_84_trigger_x_x92_symbol : Boolean;
        signal ptr_deref_84_active_x_x93_symbol : Boolean;
        signal ptr_deref_84_base_address_calculated_94_symbol : Boolean;
        signal ptr_deref_84_root_address_calculated_95_symbol : Boolean;
        signal ptr_deref_84_word_address_calculated_96_symbol : Boolean;
        signal ptr_deref_84_request_97_symbol : Boolean;
        signal ptr_deref_84_complete_108_symbol : Boolean;
        signal assign_stmt_90_active_x_x121_symbol : Boolean;
        signal assign_stmt_90_completed_x_x122_symbol : Boolean;
        signal array_obj_ref_89_trigger_x_x123_symbol : Boolean;
        signal array_obj_ref_89_active_x_x124_symbol : Boolean;
        signal array_obj_ref_89_base_address_calculated_125_symbol : Boolean;
        signal array_obj_ref_89_root_address_calculated_126_symbol : Boolean;
        signal array_obj_ref_89_base_address_resized_127_symbol : Boolean;
        signal array_obj_ref_89_base_addr_resize_128_symbol : Boolean;
        signal array_obj_ref_89_base_plus_offset_trigger_133_symbol : Boolean;
        signal array_obj_ref_89_base_plus_offset_134_symbol : Boolean;
        signal array_obj_ref_89_complete_141_symbol : Boolean;
        signal assign_stmt_94_active_x_x146_symbol : Boolean;
        signal assign_stmt_94_completed_x_x147_symbol : Boolean;
        signal ptr_deref_93_trigger_x_x148_symbol : Boolean;
        signal ptr_deref_93_active_x_x149_symbol : Boolean;
        signal ptr_deref_93_base_address_calculated_150_symbol : Boolean;
        signal simple_obj_ref_92_complete_151_symbol : Boolean;
        signal ptr_deref_93_root_address_calculated_152_symbol : Boolean;
        signal ptr_deref_93_word_address_calculated_153_symbol : Boolean;
        signal ptr_deref_93_base_address_resized_154_symbol : Boolean;
        signal ptr_deref_93_base_addr_resize_155_symbol : Boolean;
        signal ptr_deref_93_base_plus_offset_160_symbol : Boolean;
        signal ptr_deref_93_word_addrgen_165_symbol : Boolean;
        signal ptr_deref_93_request_170_symbol : Boolean;
        signal ptr_deref_93_complete_181_symbol : Boolean;
        signal assign_stmt_99_active_x_x194_symbol : Boolean;
        signal assign_stmt_99_completed_x_x195_symbol : Boolean;
        signal binary_98_active_x_x196_symbol : Boolean;
        signal binary_98_trigger_x_x197_symbol : Boolean;
        signal simple_obj_ref_97_complete_198_symbol : Boolean;
        signal binary_98_complete_199_symbol : Boolean;
        signal assign_stmt_103_active_x_x206_symbol : Boolean;
        signal assign_stmt_103_completed_x_x207_symbol : Boolean;
        signal ptr_deref_102_trigger_x_x208_symbol : Boolean;
        signal ptr_deref_102_active_x_x209_symbol : Boolean;
        signal ptr_deref_102_base_address_calculated_210_symbol : Boolean;
        signal ptr_deref_102_root_address_calculated_211_symbol : Boolean;
        signal ptr_deref_102_word_address_calculated_212_symbol : Boolean;
        signal ptr_deref_102_request_213_symbol : Boolean;
        signal ptr_deref_102_complete_224_symbol : Boolean;
        signal assign_stmt_108_active_x_x237_symbol : Boolean;
        signal assign_stmt_108_completed_x_x238_symbol : Boolean;
        signal array_obj_ref_107_trigger_x_x239_symbol : Boolean;
        signal array_obj_ref_107_active_x_x240_symbol : Boolean;
        signal array_obj_ref_107_base_address_calculated_241_symbol : Boolean;
        signal array_obj_ref_107_root_address_calculated_242_symbol : Boolean;
        signal array_obj_ref_107_base_address_resized_243_symbol : Boolean;
        signal array_obj_ref_107_base_addr_resize_244_symbol : Boolean;
        signal array_obj_ref_107_base_plus_offset_trigger_249_symbol : Boolean;
        signal array_obj_ref_107_base_plus_offset_250_symbol : Boolean;
        signal array_obj_ref_107_complete_257_symbol : Boolean;
        signal assign_stmt_112_active_x_x262_symbol : Boolean;
        signal assign_stmt_112_completed_x_x263_symbol : Boolean;
        signal simple_obj_ref_111_complete_264_symbol : Boolean;
        signal ptr_deref_110_trigger_x_x265_symbol : Boolean;
        signal ptr_deref_110_active_x_x266_symbol : Boolean;
        signal ptr_deref_110_base_address_calculated_267_symbol : Boolean;
        signal simple_obj_ref_109_complete_268_symbol : Boolean;
        signal ptr_deref_110_root_address_calculated_269_symbol : Boolean;
        signal ptr_deref_110_word_address_calculated_270_symbol : Boolean;
        signal ptr_deref_110_base_address_resized_271_symbol : Boolean;
        signal ptr_deref_110_base_addr_resize_272_symbol : Boolean;
        signal ptr_deref_110_base_plus_offset_277_symbol : Boolean;
        signal ptr_deref_110_word_addrgen_282_symbol : Boolean;
        signal ptr_deref_110_request_287_symbol : Boolean;
        signal ptr_deref_110_complete_300_symbol : Boolean;
        signal assign_stmt_116_active_x_x311_symbol : Boolean;
        signal assign_stmt_116_completed_x_x312_symbol : Boolean;
        signal ptr_deref_115_trigger_x_x313_symbol : Boolean;
        signal ptr_deref_115_active_x_x314_symbol : Boolean;
        signal ptr_deref_115_base_address_calculated_315_symbol : Boolean;
        signal ptr_deref_115_root_address_calculated_316_symbol : Boolean;
        signal ptr_deref_115_word_address_calculated_317_symbol : Boolean;
        signal ptr_deref_115_request_318_symbol : Boolean;
        signal ptr_deref_115_complete_329_symbol : Boolean;
        signal assign_stmt_120_active_x_x342_symbol : Boolean;
        signal assign_stmt_120_completed_x_x343_symbol : Boolean;
        signal type_cast_119_active_x_x344_symbol : Boolean;
        signal type_cast_119_trigger_x_x345_symbol : Boolean;
        signal simple_obj_ref_118_complete_346_symbol : Boolean;
        signal type_cast_119_complete_347_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_77_to_assign_stmt_125_45_start <= assign_stmt_77_to_assign_stmt_125_x_xentry_x_xx_x16_symbol; -- control passed to block
        Xentry_46_symbol  <= assign_stmt_77_to_assign_stmt_125_45_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/$entry
        assign_stmt_77_active_x_x48_symbol <= type_cast_76_complete_53_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_77_active_
        assign_stmt_77_completed_x_x49_symbol <= assign_stmt_77_active_x_x48_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_77_completed_
        type_cast_76_active_x_x50_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_active_ 
          signal type_cast_76_active_x_x50_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_76_active_x_x50_predecessors(0) <= type_cast_76_trigger_x_x51_symbol;
          type_cast_76_active_x_x50_predecessors(1) <= simple_obj_ref_75_complete_52_symbol;
          type_cast_76_active_x_x50_join: join -- 
            port map( -- 
              preds => type_cast_76_active_x_x50_predecessors,
              symbol_out => type_cast_76_active_x_x50_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_active_
        type_cast_76_trigger_x_x51_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_trigger_
        simple_obj_ref_75_complete_52_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_75_complete
        type_cast_76_complete_53: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete 
          signal type_cast_76_complete_53_start: Boolean;
          signal Xentry_54_symbol: Boolean;
          signal Xexit_55_symbol: Boolean;
          signal req_56_symbol : Boolean;
          signal ack_57_symbol : Boolean;
          -- 
        begin -- 
          type_cast_76_complete_53_start <= type_cast_76_active_x_x50_symbol; -- control passed to block
          Xentry_54_symbol  <= type_cast_76_complete_53_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/$entry
          req_56_symbol <= Xentry_54_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/req
          type_cast_76_inst_req_0 <= req_56_symbol; -- link to DP
          ack_57_symbol <= type_cast_76_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/ack
          Xexit_55_symbol <= ack_57_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete/$exit
          type_cast_76_complete_53_symbol <= Xexit_55_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_76_complete
        assign_stmt_81_active_x_x58_symbol <= simple_obj_ref_80_complete_60_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_81_active_
        assign_stmt_81_completed_x_x59_symbol <= ptr_deref_79_complete_79_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_81_completed_
        simple_obj_ref_80_complete_60_symbol <= assign_stmt_77_completed_x_x49_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_80_complete
        ptr_deref_79_trigger_x_x61_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_trigger_ 
          signal ptr_deref_79_trigger_x_x61_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_79_trigger_x_x61_predecessors(0) <= ptr_deref_79_word_address_calculated_65_symbol;
          ptr_deref_79_trigger_x_x61_predecessors(1) <= assign_stmt_81_active_x_x58_symbol;
          ptr_deref_79_trigger_x_x61_join: join -- 
            port map( -- 
              preds => ptr_deref_79_trigger_x_x61_predecessors,
              symbol_out => ptr_deref_79_trigger_x_x61_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_trigger_
        ptr_deref_79_active_x_x62_symbol <= ptr_deref_79_request_66_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_active_
        ptr_deref_79_base_address_calculated_63_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_base_address_calculated
        ptr_deref_79_root_address_calculated_64_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_root_address_calculated
        ptr_deref_79_word_address_calculated_65_symbol <= ptr_deref_79_root_address_calculated_64_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_word_address_calculated
        ptr_deref_79_request_66: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request 
          signal ptr_deref_79_request_66_start: Boolean;
          signal Xentry_67_symbol: Boolean;
          signal Xexit_68_symbol: Boolean;
          signal split_req_69_symbol : Boolean;
          signal split_ack_70_symbol : Boolean;
          signal word_access_71_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_79_request_66_start <= ptr_deref_79_trigger_x_x61_symbol; -- control passed to block
          Xentry_67_symbol  <= ptr_deref_79_request_66_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/$entry
          split_req_69_symbol <= Xentry_67_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/split_req
          ptr_deref_79_gather_scatter_req_0 <= split_req_69_symbol; -- link to DP
          split_ack_70_symbol <= ptr_deref_79_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/split_ack
          word_access_71: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access 
            signal word_access_71_start: Boolean;
            signal Xentry_72_symbol: Boolean;
            signal Xexit_73_symbol: Boolean;
            signal word_access_0_74_symbol : Boolean;
            -- 
          begin -- 
            word_access_71_start <= split_ack_70_symbol; -- control passed to block
            Xentry_72_symbol  <= word_access_71_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/$entry
            word_access_0_74: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0 
              signal word_access_0_74_start: Boolean;
              signal Xentry_75_symbol: Boolean;
              signal Xexit_76_symbol: Boolean;
              signal rr_77_symbol : Boolean;
              signal ra_78_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_74_start <= Xentry_72_symbol; -- control passed to block
              Xentry_75_symbol  <= word_access_0_74_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/$entry
              rr_77_symbol <= Xentry_75_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/rr
              ptr_deref_79_store_0_req_0 <= rr_77_symbol; -- link to DP
              ra_78_symbol <= ptr_deref_79_store_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/ra
              Xexit_76_symbol <= ra_78_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0/$exit
              word_access_0_74_symbol <= Xexit_76_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/word_access_0
            Xexit_73_symbol <= word_access_0_74_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access/$exit
            word_access_71_symbol <= Xexit_73_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/word_access
          Xexit_68_symbol <= word_access_71_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request/$exit
          ptr_deref_79_request_66_symbol <= Xexit_68_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_request
        ptr_deref_79_complete_79: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete 
          signal ptr_deref_79_complete_79_start: Boolean;
          signal Xentry_80_symbol: Boolean;
          signal Xexit_81_symbol: Boolean;
          signal word_access_82_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_79_complete_79_start <= ptr_deref_79_active_x_x62_symbol; -- control passed to block
          Xentry_80_symbol  <= ptr_deref_79_complete_79_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/$entry
          word_access_82: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access 
            signal word_access_82_start: Boolean;
            signal Xentry_83_symbol: Boolean;
            signal Xexit_84_symbol: Boolean;
            signal word_access_0_85_symbol : Boolean;
            -- 
          begin -- 
            word_access_82_start <= Xentry_80_symbol; -- control passed to block
            Xentry_83_symbol  <= word_access_82_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/$entry
            word_access_0_85: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0 
              signal word_access_0_85_start: Boolean;
              signal Xentry_86_symbol: Boolean;
              signal Xexit_87_symbol: Boolean;
              signal cr_88_symbol : Boolean;
              signal ca_89_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_85_start <= Xentry_83_symbol; -- control passed to block
              Xentry_86_symbol  <= word_access_0_85_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/$entry
              cr_88_symbol <= Xentry_86_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/cr
              ptr_deref_79_store_0_req_1 <= cr_88_symbol; -- link to DP
              ca_89_symbol <= ptr_deref_79_store_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/ca
              Xexit_87_symbol <= ca_89_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0/$exit
              word_access_0_85_symbol <= Xexit_87_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/word_access_0
            Xexit_84_symbol <= word_access_0_85_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access/$exit
            word_access_82_symbol <= Xexit_84_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/word_access
          Xexit_81_symbol <= word_access_82_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete/$exit
          ptr_deref_79_complete_79_symbol <= Xexit_81_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_79_complete
        assign_stmt_85_active_x_x90_symbol <= ptr_deref_84_complete_108_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_85_active_
        assign_stmt_85_completed_x_x91_symbol <= assign_stmt_85_active_x_x90_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_85_completed_
        ptr_deref_84_trigger_x_x92_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_trigger_ 
          signal ptr_deref_84_trigger_x_x92_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_84_trigger_x_x92_predecessors(0) <= ptr_deref_84_word_address_calculated_96_symbol;
          ptr_deref_84_trigger_x_x92_predecessors(1) <= ptr_deref_79_active_x_x62_symbol;
          ptr_deref_84_trigger_x_x92_join: join -- 
            port map( -- 
              preds => ptr_deref_84_trigger_x_x92_predecessors,
              symbol_out => ptr_deref_84_trigger_x_x92_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_trigger_
        ptr_deref_84_active_x_x93_symbol <= ptr_deref_84_request_97_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_active_
        ptr_deref_84_base_address_calculated_94_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_base_address_calculated
        ptr_deref_84_root_address_calculated_95_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_root_address_calculated
        ptr_deref_84_word_address_calculated_96_symbol <= ptr_deref_84_root_address_calculated_95_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_word_address_calculated
        ptr_deref_84_request_97: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request 
          signal ptr_deref_84_request_97_start: Boolean;
          signal Xentry_98_symbol: Boolean;
          signal Xexit_99_symbol: Boolean;
          signal word_access_100_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_84_request_97_start <= ptr_deref_84_trigger_x_x92_symbol; -- control passed to block
          Xentry_98_symbol  <= ptr_deref_84_request_97_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/$entry
          word_access_100: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access 
            signal word_access_100_start: Boolean;
            signal Xentry_101_symbol: Boolean;
            signal Xexit_102_symbol: Boolean;
            signal word_access_0_103_symbol : Boolean;
            -- 
          begin -- 
            word_access_100_start <= Xentry_98_symbol; -- control passed to block
            Xentry_101_symbol  <= word_access_100_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/$entry
            word_access_0_103: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0 
              signal word_access_0_103_start: Boolean;
              signal Xentry_104_symbol: Boolean;
              signal Xexit_105_symbol: Boolean;
              signal rr_106_symbol : Boolean;
              signal ra_107_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_103_start <= Xentry_101_symbol; -- control passed to block
              Xentry_104_symbol  <= word_access_0_103_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/$entry
              rr_106_symbol <= Xentry_104_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/rr
              ptr_deref_84_load_0_req_0 <= rr_106_symbol; -- link to DP
              ra_107_symbol <= ptr_deref_84_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/ra
              Xexit_105_symbol <= ra_107_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0/$exit
              word_access_0_103_symbol <= Xexit_105_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/word_access_0
            Xexit_102_symbol <= word_access_0_103_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access/$exit
            word_access_100_symbol <= Xexit_102_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/word_access
          Xexit_99_symbol <= word_access_100_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request/$exit
          ptr_deref_84_request_97_symbol <= Xexit_99_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_request
        ptr_deref_84_complete_108: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete 
          signal ptr_deref_84_complete_108_start: Boolean;
          signal Xentry_109_symbol: Boolean;
          signal Xexit_110_symbol: Boolean;
          signal word_access_111_symbol : Boolean;
          signal merge_req_119_symbol : Boolean;
          signal merge_ack_120_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_84_complete_108_start <= ptr_deref_84_active_x_x93_symbol; -- control passed to block
          Xentry_109_symbol  <= ptr_deref_84_complete_108_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/$entry
          word_access_111: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access 
            signal word_access_111_start: Boolean;
            signal Xentry_112_symbol: Boolean;
            signal Xexit_113_symbol: Boolean;
            signal word_access_0_114_symbol : Boolean;
            -- 
          begin -- 
            word_access_111_start <= Xentry_109_symbol; -- control passed to block
            Xentry_112_symbol  <= word_access_111_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/$entry
            word_access_0_114: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0 
              signal word_access_0_114_start: Boolean;
              signal Xentry_115_symbol: Boolean;
              signal Xexit_116_symbol: Boolean;
              signal cr_117_symbol : Boolean;
              signal ca_118_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_114_start <= Xentry_112_symbol; -- control passed to block
              Xentry_115_symbol  <= word_access_0_114_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/$entry
              cr_117_symbol <= Xentry_115_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/cr
              ptr_deref_84_load_0_req_1 <= cr_117_symbol; -- link to DP
              ca_118_symbol <= ptr_deref_84_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/ca
              Xexit_116_symbol <= ca_118_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0/$exit
              word_access_0_114_symbol <= Xexit_116_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/word_access_0
            Xexit_113_symbol <= word_access_0_114_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access/$exit
            word_access_111_symbol <= Xexit_113_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/word_access
          merge_req_119_symbol <= word_access_111_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/merge_req
          ptr_deref_84_gather_scatter_req_0 <= merge_req_119_symbol; -- link to DP
          merge_ack_120_symbol <= ptr_deref_84_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/merge_ack
          Xexit_110_symbol <= merge_ack_120_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete/$exit
          ptr_deref_84_complete_108_symbol <= Xexit_110_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_84_complete
        assign_stmt_90_active_x_x121_symbol <= array_obj_ref_89_complete_141_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_90_active_
        assign_stmt_90_completed_x_x122_symbol <= assign_stmt_90_active_x_x121_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_90_completed_
        array_obj_ref_89_trigger_x_x123_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_trigger_
        array_obj_ref_89_active_x_x124_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_active_ 
          signal array_obj_ref_89_active_x_x124_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_89_active_x_x124_predecessors(0) <= array_obj_ref_89_trigger_x_x123_symbol;
          array_obj_ref_89_active_x_x124_predecessors(1) <= array_obj_ref_89_root_address_calculated_126_symbol;
          array_obj_ref_89_active_x_x124_join: join -- 
            port map( -- 
              preds => array_obj_ref_89_active_x_x124_predecessors,
              symbol_out => array_obj_ref_89_active_x_x124_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_active_
        array_obj_ref_89_base_address_calculated_125_symbol <= assign_stmt_85_completed_x_x91_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_address_calculated
        array_obj_ref_89_root_address_calculated_126_symbol <= array_obj_ref_89_base_plus_offset_134_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_root_address_calculated
        array_obj_ref_89_base_address_resized_127_symbol <= array_obj_ref_89_base_addr_resize_128_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_address_resized
        array_obj_ref_89_base_addr_resize_128: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize 
          signal array_obj_ref_89_base_addr_resize_128_start: Boolean;
          signal Xentry_129_symbol: Boolean;
          signal Xexit_130_symbol: Boolean;
          signal base_resize_req_131_symbol : Boolean;
          signal base_resize_ack_132_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_89_base_addr_resize_128_start <= array_obj_ref_89_base_address_calculated_125_symbol; -- control passed to block
          Xentry_129_symbol  <= array_obj_ref_89_base_addr_resize_128_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/$entry
          base_resize_req_131_symbol <= Xentry_129_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/base_resize_req
          array_obj_ref_89_base_resize_req_0 <= base_resize_req_131_symbol; -- link to DP
          base_resize_ack_132_symbol <= array_obj_ref_89_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/base_resize_ack
          Xexit_130_symbol <= base_resize_ack_132_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize/$exit
          array_obj_ref_89_base_addr_resize_128_symbol <= Xexit_130_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_addr_resize
        array_obj_ref_89_base_plus_offset_trigger_133_symbol <= array_obj_ref_89_base_address_resized_127_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset_trigger
        array_obj_ref_89_base_plus_offset_134: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset 
          signal array_obj_ref_89_base_plus_offset_134_start: Boolean;
          signal Xentry_135_symbol: Boolean;
          signal Xexit_136_symbol: Boolean;
          signal plus_base_rr_137_symbol : Boolean;
          signal plus_base_ra_138_symbol : Boolean;
          signal plus_base_cr_139_symbol : Boolean;
          signal plus_base_ca_140_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_89_base_plus_offset_134_start <= array_obj_ref_89_base_plus_offset_trigger_133_symbol; -- control passed to block
          Xentry_135_symbol  <= array_obj_ref_89_base_plus_offset_134_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/$entry
          plus_base_rr_137_symbol <= Xentry_135_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_rr
          array_obj_ref_89_root_address_inst_req_0 <= plus_base_rr_137_symbol; -- link to DP
          plus_base_ra_138_symbol <= array_obj_ref_89_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_ra
          plus_base_cr_139_symbol <= plus_base_ra_138_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_cr
          array_obj_ref_89_root_address_inst_req_1 <= plus_base_cr_139_symbol; -- link to DP
          plus_base_ca_140_symbol <= array_obj_ref_89_root_address_inst_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/plus_base_ca
          Xexit_136_symbol <= plus_base_ca_140_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset/$exit
          array_obj_ref_89_base_plus_offset_134_symbol <= Xexit_136_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_base_plus_offset
        array_obj_ref_89_complete_141: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete 
          signal array_obj_ref_89_complete_141_start: Boolean;
          signal Xentry_142_symbol: Boolean;
          signal Xexit_143_symbol: Boolean;
          signal final_reg_req_144_symbol : Boolean;
          signal final_reg_ack_145_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_89_complete_141_start <= array_obj_ref_89_active_x_x124_symbol; -- control passed to block
          Xentry_142_symbol  <= array_obj_ref_89_complete_141_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/$entry
          final_reg_req_144_symbol <= Xentry_142_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/final_reg_req
          array_obj_ref_89_final_reg_req_0 <= final_reg_req_144_symbol; -- link to DP
          final_reg_ack_145_symbol <= array_obj_ref_89_final_reg_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/final_reg_ack
          Xexit_143_symbol <= final_reg_ack_145_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete/$exit
          array_obj_ref_89_complete_141_symbol <= Xexit_143_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_89_complete
        assign_stmt_94_active_x_x146_symbol <= ptr_deref_93_complete_181_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_94_active_
        assign_stmt_94_completed_x_x147_symbol <= assign_stmt_94_active_x_x146_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_94_completed_
        ptr_deref_93_trigger_x_x148_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_trigger_ 
          signal ptr_deref_93_trigger_x_x148_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_93_trigger_x_x148_predecessors(0) <= ptr_deref_93_word_address_calculated_153_symbol;
          ptr_deref_93_trigger_x_x148_predecessors(1) <= ptr_deref_93_base_address_calculated_150_symbol;
          ptr_deref_93_trigger_x_x148_join: join -- 
            port map( -- 
              preds => ptr_deref_93_trigger_x_x148_predecessors,
              symbol_out => ptr_deref_93_trigger_x_x148_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_trigger_
        ptr_deref_93_active_x_x149_symbol <= ptr_deref_93_request_170_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_active_
        ptr_deref_93_base_address_calculated_150_symbol <= simple_obj_ref_92_complete_151_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_address_calculated
        simple_obj_ref_92_complete_151_symbol <= assign_stmt_90_completed_x_x122_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_92_complete
        ptr_deref_93_root_address_calculated_152_symbol <= ptr_deref_93_base_plus_offset_160_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_root_address_calculated
        ptr_deref_93_word_address_calculated_153_symbol <= ptr_deref_93_word_addrgen_165_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_address_calculated
        ptr_deref_93_base_address_resized_154_symbol <= ptr_deref_93_base_addr_resize_155_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_address_resized
        ptr_deref_93_base_addr_resize_155: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize 
          signal ptr_deref_93_base_addr_resize_155_start: Boolean;
          signal Xentry_156_symbol: Boolean;
          signal Xexit_157_symbol: Boolean;
          signal base_resize_req_158_symbol : Boolean;
          signal base_resize_ack_159_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_base_addr_resize_155_start <= ptr_deref_93_base_address_calculated_150_symbol; -- control passed to block
          Xentry_156_symbol  <= ptr_deref_93_base_addr_resize_155_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/$entry
          base_resize_req_158_symbol <= Xentry_156_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/base_resize_req
          ptr_deref_93_base_resize_req_0 <= base_resize_req_158_symbol; -- link to DP
          base_resize_ack_159_symbol <= ptr_deref_93_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/base_resize_ack
          Xexit_157_symbol <= base_resize_ack_159_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize/$exit
          ptr_deref_93_base_addr_resize_155_symbol <= Xexit_157_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_addr_resize
        ptr_deref_93_base_plus_offset_160: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset 
          signal ptr_deref_93_base_plus_offset_160_start: Boolean;
          signal Xentry_161_symbol: Boolean;
          signal Xexit_162_symbol: Boolean;
          signal sum_rename_req_163_symbol : Boolean;
          signal sum_rename_ack_164_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_base_plus_offset_160_start <= ptr_deref_93_base_address_resized_154_symbol; -- control passed to block
          Xentry_161_symbol  <= ptr_deref_93_base_plus_offset_160_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/$entry
          sum_rename_req_163_symbol <= Xentry_161_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/sum_rename_req
          ptr_deref_93_root_address_inst_req_0 <= sum_rename_req_163_symbol; -- link to DP
          sum_rename_ack_164_symbol <= ptr_deref_93_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/sum_rename_ack
          Xexit_162_symbol <= sum_rename_ack_164_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset/$exit
          ptr_deref_93_base_plus_offset_160_symbol <= Xexit_162_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_base_plus_offset
        ptr_deref_93_word_addrgen_165: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen 
          signal ptr_deref_93_word_addrgen_165_start: Boolean;
          signal Xentry_166_symbol: Boolean;
          signal Xexit_167_symbol: Boolean;
          signal root_rename_req_168_symbol : Boolean;
          signal root_rename_ack_169_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_word_addrgen_165_start <= ptr_deref_93_root_address_calculated_152_symbol; -- control passed to block
          Xentry_166_symbol  <= ptr_deref_93_word_addrgen_165_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/$entry
          root_rename_req_168_symbol <= Xentry_166_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/root_rename_req
          ptr_deref_93_addr_0_req_0 <= root_rename_req_168_symbol; -- link to DP
          root_rename_ack_169_symbol <= ptr_deref_93_addr_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/root_rename_ack
          Xexit_167_symbol <= root_rename_ack_169_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen/$exit
          ptr_deref_93_word_addrgen_165_symbol <= Xexit_167_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_word_addrgen
        ptr_deref_93_request_170: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request 
          signal ptr_deref_93_request_170_start: Boolean;
          signal Xentry_171_symbol: Boolean;
          signal Xexit_172_symbol: Boolean;
          signal word_access_173_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_request_170_start <= ptr_deref_93_trigger_x_x148_symbol; -- control passed to block
          Xentry_171_symbol  <= ptr_deref_93_request_170_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/$entry
          word_access_173: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access 
            signal word_access_173_start: Boolean;
            signal Xentry_174_symbol: Boolean;
            signal Xexit_175_symbol: Boolean;
            signal word_access_0_176_symbol : Boolean;
            -- 
          begin -- 
            word_access_173_start <= Xentry_171_symbol; -- control passed to block
            Xentry_174_symbol  <= word_access_173_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/$entry
            word_access_0_176: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0 
              signal word_access_0_176_start: Boolean;
              signal Xentry_177_symbol: Boolean;
              signal Xexit_178_symbol: Boolean;
              signal rr_179_symbol : Boolean;
              signal ra_180_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_176_start <= Xentry_174_symbol; -- control passed to block
              Xentry_177_symbol  <= word_access_0_176_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/$entry
              rr_179_symbol <= Xentry_177_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/rr
              ptr_deref_93_load_0_req_0 <= rr_179_symbol; -- link to DP
              ra_180_symbol <= ptr_deref_93_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/ra
              Xexit_178_symbol <= ra_180_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0/$exit
              word_access_0_176_symbol <= Xexit_178_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/word_access_0
            Xexit_175_symbol <= word_access_0_176_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access/$exit
            word_access_173_symbol <= Xexit_175_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/word_access
          Xexit_172_symbol <= word_access_173_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request/$exit
          ptr_deref_93_request_170_symbol <= Xexit_172_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_request
        ptr_deref_93_complete_181: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete 
          signal ptr_deref_93_complete_181_start: Boolean;
          signal Xentry_182_symbol: Boolean;
          signal Xexit_183_symbol: Boolean;
          signal word_access_184_symbol : Boolean;
          signal merge_req_192_symbol : Boolean;
          signal merge_ack_193_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_93_complete_181_start <= ptr_deref_93_active_x_x149_symbol; -- control passed to block
          Xentry_182_symbol  <= ptr_deref_93_complete_181_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/$entry
          word_access_184: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access 
            signal word_access_184_start: Boolean;
            signal Xentry_185_symbol: Boolean;
            signal Xexit_186_symbol: Boolean;
            signal word_access_0_187_symbol : Boolean;
            -- 
          begin -- 
            word_access_184_start <= Xentry_182_symbol; -- control passed to block
            Xentry_185_symbol  <= word_access_184_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/$entry
            word_access_0_187: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0 
              signal word_access_0_187_start: Boolean;
              signal Xentry_188_symbol: Boolean;
              signal Xexit_189_symbol: Boolean;
              signal cr_190_symbol : Boolean;
              signal ca_191_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_187_start <= Xentry_185_symbol; -- control passed to block
              Xentry_188_symbol  <= word_access_0_187_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/$entry
              cr_190_symbol <= Xentry_188_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/cr
              ptr_deref_93_load_0_req_1 <= cr_190_symbol; -- link to DP
              ca_191_symbol <= ptr_deref_93_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/ca
              Xexit_189_symbol <= ca_191_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0/$exit
              word_access_0_187_symbol <= Xexit_189_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/word_access_0
            Xexit_186_symbol <= word_access_0_187_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access/$exit
            word_access_184_symbol <= Xexit_186_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/word_access
          merge_req_192_symbol <= word_access_184_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/merge_req
          ptr_deref_93_gather_scatter_req_0 <= merge_req_192_symbol; -- link to DP
          merge_ack_193_symbol <= ptr_deref_93_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/merge_ack
          Xexit_183_symbol <= merge_ack_193_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete/$exit
          ptr_deref_93_complete_181_symbol <= Xexit_183_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_93_complete
        assign_stmt_99_active_x_x194_symbol <= binary_98_complete_199_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_99_active_
        assign_stmt_99_completed_x_x195_symbol <= assign_stmt_99_active_x_x194_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_99_completed_
        binary_98_active_x_x196_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_active_ 
          signal binary_98_active_x_x196_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_98_active_x_x196_predecessors(0) <= binary_98_trigger_x_x197_symbol;
          binary_98_active_x_x196_predecessors(1) <= simple_obj_ref_97_complete_198_symbol;
          binary_98_active_x_x196_join: join -- 
            port map( -- 
              preds => binary_98_active_x_x196_predecessors,
              symbol_out => binary_98_active_x_x196_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_active_
        binary_98_trigger_x_x197_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_trigger_
        simple_obj_ref_97_complete_198_symbol <= assign_stmt_94_completed_x_x147_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_97_complete
        binary_98_complete_199: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete 
          signal binary_98_complete_199_start: Boolean;
          signal Xentry_200_symbol: Boolean;
          signal Xexit_201_symbol: Boolean;
          signal rr_202_symbol : Boolean;
          signal ra_203_symbol : Boolean;
          signal cr_204_symbol : Boolean;
          signal ca_205_symbol : Boolean;
          -- 
        begin -- 
          binary_98_complete_199_start <= binary_98_active_x_x196_symbol; -- control passed to block
          Xentry_200_symbol  <= binary_98_complete_199_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/$entry
          rr_202_symbol <= Xentry_200_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/rr
          binary_98_inst_req_0 <= rr_202_symbol; -- link to DP
          ra_203_symbol <= binary_98_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/ra
          cr_204_symbol <= ra_203_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/cr
          binary_98_inst_req_1 <= cr_204_symbol; -- link to DP
          ca_205_symbol <= binary_98_inst_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/ca
          Xexit_201_symbol <= ca_205_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete/$exit
          binary_98_complete_199_symbol <= Xexit_201_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/binary_98_complete
        assign_stmt_103_active_x_x206_symbol <= ptr_deref_102_complete_224_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_103_active_
        assign_stmt_103_completed_x_x207_symbol <= assign_stmt_103_active_x_x206_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_103_completed_
        ptr_deref_102_trigger_x_x208_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_trigger_ 
          signal ptr_deref_102_trigger_x_x208_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_102_trigger_x_x208_predecessors(0) <= ptr_deref_102_word_address_calculated_212_symbol;
          ptr_deref_102_trigger_x_x208_predecessors(1) <= ptr_deref_79_active_x_x62_symbol;
          ptr_deref_102_trigger_x_x208_join: join -- 
            port map( -- 
              preds => ptr_deref_102_trigger_x_x208_predecessors,
              symbol_out => ptr_deref_102_trigger_x_x208_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_trigger_
        ptr_deref_102_active_x_x209_symbol <= ptr_deref_102_request_213_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_active_
        ptr_deref_102_base_address_calculated_210_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_base_address_calculated
        ptr_deref_102_root_address_calculated_211_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_root_address_calculated
        ptr_deref_102_word_address_calculated_212_symbol <= ptr_deref_102_root_address_calculated_211_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_word_address_calculated
        ptr_deref_102_request_213: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request 
          signal ptr_deref_102_request_213_start: Boolean;
          signal Xentry_214_symbol: Boolean;
          signal Xexit_215_symbol: Boolean;
          signal word_access_216_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_102_request_213_start <= ptr_deref_102_trigger_x_x208_symbol; -- control passed to block
          Xentry_214_symbol  <= ptr_deref_102_request_213_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/$entry
          word_access_216: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access 
            signal word_access_216_start: Boolean;
            signal Xentry_217_symbol: Boolean;
            signal Xexit_218_symbol: Boolean;
            signal word_access_0_219_symbol : Boolean;
            -- 
          begin -- 
            word_access_216_start <= Xentry_214_symbol; -- control passed to block
            Xentry_217_symbol  <= word_access_216_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/$entry
            word_access_0_219: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0 
              signal word_access_0_219_start: Boolean;
              signal Xentry_220_symbol: Boolean;
              signal Xexit_221_symbol: Boolean;
              signal rr_222_symbol : Boolean;
              signal ra_223_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_219_start <= Xentry_217_symbol; -- control passed to block
              Xentry_220_symbol  <= word_access_0_219_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/$entry
              rr_222_symbol <= Xentry_220_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/rr
              ptr_deref_102_load_0_req_0 <= rr_222_symbol; -- link to DP
              ra_223_symbol <= ptr_deref_102_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/ra
              Xexit_221_symbol <= ra_223_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0/$exit
              word_access_0_219_symbol <= Xexit_221_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/word_access_0
            Xexit_218_symbol <= word_access_0_219_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access/$exit
            word_access_216_symbol <= Xexit_218_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/word_access
          Xexit_215_symbol <= word_access_216_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request/$exit
          ptr_deref_102_request_213_symbol <= Xexit_215_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_request
        ptr_deref_102_complete_224: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete 
          signal ptr_deref_102_complete_224_start: Boolean;
          signal Xentry_225_symbol: Boolean;
          signal Xexit_226_symbol: Boolean;
          signal word_access_227_symbol : Boolean;
          signal merge_req_235_symbol : Boolean;
          signal merge_ack_236_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_102_complete_224_start <= ptr_deref_102_active_x_x209_symbol; -- control passed to block
          Xentry_225_symbol  <= ptr_deref_102_complete_224_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/$entry
          word_access_227: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access 
            signal word_access_227_start: Boolean;
            signal Xentry_228_symbol: Boolean;
            signal Xexit_229_symbol: Boolean;
            signal word_access_0_230_symbol : Boolean;
            -- 
          begin -- 
            word_access_227_start <= Xentry_225_symbol; -- control passed to block
            Xentry_228_symbol  <= word_access_227_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/$entry
            word_access_0_230: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0 
              signal word_access_0_230_start: Boolean;
              signal Xentry_231_symbol: Boolean;
              signal Xexit_232_symbol: Boolean;
              signal cr_233_symbol : Boolean;
              signal ca_234_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_230_start <= Xentry_228_symbol; -- control passed to block
              Xentry_231_symbol  <= word_access_0_230_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/$entry
              cr_233_symbol <= Xentry_231_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/cr
              ptr_deref_102_load_0_req_1 <= cr_233_symbol; -- link to DP
              ca_234_symbol <= ptr_deref_102_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/ca
              Xexit_232_symbol <= ca_234_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0/$exit
              word_access_0_230_symbol <= Xexit_232_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/word_access_0
            Xexit_229_symbol <= word_access_0_230_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access/$exit
            word_access_227_symbol <= Xexit_229_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/word_access
          merge_req_235_symbol <= word_access_227_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/merge_req
          ptr_deref_102_gather_scatter_req_0 <= merge_req_235_symbol; -- link to DP
          merge_ack_236_symbol <= ptr_deref_102_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/merge_ack
          Xexit_226_symbol <= merge_ack_236_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete/$exit
          ptr_deref_102_complete_224_symbol <= Xexit_226_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_102_complete
        assign_stmt_108_active_x_x237_symbol <= array_obj_ref_107_complete_257_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_108_active_
        assign_stmt_108_completed_x_x238_symbol <= assign_stmt_108_active_x_x237_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_108_completed_
        array_obj_ref_107_trigger_x_x239_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_trigger_
        array_obj_ref_107_active_x_x240_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_active_ 
          signal array_obj_ref_107_active_x_x240_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_107_active_x_x240_predecessors(0) <= array_obj_ref_107_trigger_x_x239_symbol;
          array_obj_ref_107_active_x_x240_predecessors(1) <= array_obj_ref_107_root_address_calculated_242_symbol;
          array_obj_ref_107_active_x_x240_join: join -- 
            port map( -- 
              preds => array_obj_ref_107_active_x_x240_predecessors,
              symbol_out => array_obj_ref_107_active_x_x240_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_active_
        array_obj_ref_107_base_address_calculated_241_symbol <= assign_stmt_103_completed_x_x207_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_address_calculated
        array_obj_ref_107_root_address_calculated_242_symbol <= array_obj_ref_107_base_plus_offset_250_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_root_address_calculated
        array_obj_ref_107_base_address_resized_243_symbol <= array_obj_ref_107_base_addr_resize_244_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_address_resized
        array_obj_ref_107_base_addr_resize_244: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize 
          signal array_obj_ref_107_base_addr_resize_244_start: Boolean;
          signal Xentry_245_symbol: Boolean;
          signal Xexit_246_symbol: Boolean;
          signal base_resize_req_247_symbol : Boolean;
          signal base_resize_ack_248_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_107_base_addr_resize_244_start <= array_obj_ref_107_base_address_calculated_241_symbol; -- control passed to block
          Xentry_245_symbol  <= array_obj_ref_107_base_addr_resize_244_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/$entry
          base_resize_req_247_symbol <= Xentry_245_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/base_resize_req
          array_obj_ref_107_base_resize_req_0 <= base_resize_req_247_symbol; -- link to DP
          base_resize_ack_248_symbol <= array_obj_ref_107_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/base_resize_ack
          Xexit_246_symbol <= base_resize_ack_248_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize/$exit
          array_obj_ref_107_base_addr_resize_244_symbol <= Xexit_246_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_addr_resize
        array_obj_ref_107_base_plus_offset_trigger_249_symbol <= array_obj_ref_107_base_address_resized_243_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset_trigger
        array_obj_ref_107_base_plus_offset_250: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset 
          signal array_obj_ref_107_base_plus_offset_250_start: Boolean;
          signal Xentry_251_symbol: Boolean;
          signal Xexit_252_symbol: Boolean;
          signal plus_base_rr_253_symbol : Boolean;
          signal plus_base_ra_254_symbol : Boolean;
          signal plus_base_cr_255_symbol : Boolean;
          signal plus_base_ca_256_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_107_base_plus_offset_250_start <= array_obj_ref_107_base_plus_offset_trigger_249_symbol; -- control passed to block
          Xentry_251_symbol  <= array_obj_ref_107_base_plus_offset_250_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/$entry
          plus_base_rr_253_symbol <= Xentry_251_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_rr
          array_obj_ref_107_root_address_inst_req_0 <= plus_base_rr_253_symbol; -- link to DP
          plus_base_ra_254_symbol <= array_obj_ref_107_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_ra
          plus_base_cr_255_symbol <= plus_base_ra_254_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_cr
          array_obj_ref_107_root_address_inst_req_1 <= plus_base_cr_255_symbol; -- link to DP
          plus_base_ca_256_symbol <= array_obj_ref_107_root_address_inst_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/plus_base_ca
          Xexit_252_symbol <= plus_base_ca_256_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset/$exit
          array_obj_ref_107_base_plus_offset_250_symbol <= Xexit_252_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_base_plus_offset
        array_obj_ref_107_complete_257: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete 
          signal array_obj_ref_107_complete_257_start: Boolean;
          signal Xentry_258_symbol: Boolean;
          signal Xexit_259_symbol: Boolean;
          signal final_reg_req_260_symbol : Boolean;
          signal final_reg_ack_261_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_107_complete_257_start <= array_obj_ref_107_active_x_x240_symbol; -- control passed to block
          Xentry_258_symbol  <= array_obj_ref_107_complete_257_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/$entry
          final_reg_req_260_symbol <= Xentry_258_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/final_reg_req
          array_obj_ref_107_final_reg_req_0 <= final_reg_req_260_symbol; -- link to DP
          final_reg_ack_261_symbol <= array_obj_ref_107_final_reg_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/final_reg_ack
          Xexit_259_symbol <= final_reg_ack_261_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete/$exit
          array_obj_ref_107_complete_257_symbol <= Xexit_259_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/array_obj_ref_107_complete
        assign_stmt_112_active_x_x262_symbol <= simple_obj_ref_111_complete_264_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_112_active_
        assign_stmt_112_completed_x_x263_symbol <= ptr_deref_110_complete_300_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_112_completed_
        simple_obj_ref_111_complete_264_symbol <= assign_stmt_99_completed_x_x195_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_111_complete
        ptr_deref_110_trigger_x_x265_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_trigger_ 
          signal ptr_deref_110_trigger_x_x265_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          ptr_deref_110_trigger_x_x265_predecessors(0) <= ptr_deref_110_word_address_calculated_270_symbol;
          ptr_deref_110_trigger_x_x265_predecessors(1) <= ptr_deref_110_base_address_calculated_267_symbol;
          ptr_deref_110_trigger_x_x265_predecessors(2) <= assign_stmt_112_active_x_x262_symbol;
          ptr_deref_110_trigger_x_x265_predecessors(3) <= ptr_deref_93_active_x_x149_symbol;
          ptr_deref_110_trigger_x_x265_join: join -- 
            port map( -- 
              preds => ptr_deref_110_trigger_x_x265_predecessors,
              symbol_out => ptr_deref_110_trigger_x_x265_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_trigger_
        ptr_deref_110_active_x_x266_symbol <= ptr_deref_110_request_287_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_active_
        ptr_deref_110_base_address_calculated_267_symbol <= simple_obj_ref_109_complete_268_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_address_calculated
        simple_obj_ref_109_complete_268_symbol <= assign_stmt_108_completed_x_x238_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_109_complete
        ptr_deref_110_root_address_calculated_269_symbol <= ptr_deref_110_base_plus_offset_277_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_root_address_calculated
        ptr_deref_110_word_address_calculated_270_symbol <= ptr_deref_110_word_addrgen_282_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_address_calculated
        ptr_deref_110_base_address_resized_271_symbol <= ptr_deref_110_base_addr_resize_272_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_address_resized
        ptr_deref_110_base_addr_resize_272: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize 
          signal ptr_deref_110_base_addr_resize_272_start: Boolean;
          signal Xentry_273_symbol: Boolean;
          signal Xexit_274_symbol: Boolean;
          signal base_resize_req_275_symbol : Boolean;
          signal base_resize_ack_276_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_base_addr_resize_272_start <= ptr_deref_110_base_address_calculated_267_symbol; -- control passed to block
          Xentry_273_symbol  <= ptr_deref_110_base_addr_resize_272_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/$entry
          base_resize_req_275_symbol <= Xentry_273_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/base_resize_req
          ptr_deref_110_base_resize_req_0 <= base_resize_req_275_symbol; -- link to DP
          base_resize_ack_276_symbol <= ptr_deref_110_base_resize_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/base_resize_ack
          Xexit_274_symbol <= base_resize_ack_276_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize/$exit
          ptr_deref_110_base_addr_resize_272_symbol <= Xexit_274_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_addr_resize
        ptr_deref_110_base_plus_offset_277: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset 
          signal ptr_deref_110_base_plus_offset_277_start: Boolean;
          signal Xentry_278_symbol: Boolean;
          signal Xexit_279_symbol: Boolean;
          signal sum_rename_req_280_symbol : Boolean;
          signal sum_rename_ack_281_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_base_plus_offset_277_start <= ptr_deref_110_base_address_resized_271_symbol; -- control passed to block
          Xentry_278_symbol  <= ptr_deref_110_base_plus_offset_277_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/$entry
          sum_rename_req_280_symbol <= Xentry_278_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/sum_rename_req
          ptr_deref_110_root_address_inst_req_0 <= sum_rename_req_280_symbol; -- link to DP
          sum_rename_ack_281_symbol <= ptr_deref_110_root_address_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/sum_rename_ack
          Xexit_279_symbol <= sum_rename_ack_281_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset/$exit
          ptr_deref_110_base_plus_offset_277_symbol <= Xexit_279_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_base_plus_offset
        ptr_deref_110_word_addrgen_282: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen 
          signal ptr_deref_110_word_addrgen_282_start: Boolean;
          signal Xentry_283_symbol: Boolean;
          signal Xexit_284_symbol: Boolean;
          signal root_rename_req_285_symbol : Boolean;
          signal root_rename_ack_286_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_word_addrgen_282_start <= ptr_deref_110_root_address_calculated_269_symbol; -- control passed to block
          Xentry_283_symbol  <= ptr_deref_110_word_addrgen_282_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/$entry
          root_rename_req_285_symbol <= Xentry_283_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/root_rename_req
          ptr_deref_110_addr_0_req_0 <= root_rename_req_285_symbol; -- link to DP
          root_rename_ack_286_symbol <= ptr_deref_110_addr_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/root_rename_ack
          Xexit_284_symbol <= root_rename_ack_286_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen/$exit
          ptr_deref_110_word_addrgen_282_symbol <= Xexit_284_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_word_addrgen
        ptr_deref_110_request_287: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request 
          signal ptr_deref_110_request_287_start: Boolean;
          signal Xentry_288_symbol: Boolean;
          signal Xexit_289_symbol: Boolean;
          signal split_req_290_symbol : Boolean;
          signal split_ack_291_symbol : Boolean;
          signal word_access_292_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_request_287_start <= ptr_deref_110_trigger_x_x265_symbol; -- control passed to block
          Xentry_288_symbol  <= ptr_deref_110_request_287_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/$entry
          split_req_290_symbol <= Xentry_288_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/split_req
          ptr_deref_110_gather_scatter_req_0 <= split_req_290_symbol; -- link to DP
          split_ack_291_symbol <= ptr_deref_110_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/split_ack
          word_access_292: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access 
            signal word_access_292_start: Boolean;
            signal Xentry_293_symbol: Boolean;
            signal Xexit_294_symbol: Boolean;
            signal word_access_0_295_symbol : Boolean;
            -- 
          begin -- 
            word_access_292_start <= split_ack_291_symbol; -- control passed to block
            Xentry_293_symbol  <= word_access_292_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/$entry
            word_access_0_295: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0 
              signal word_access_0_295_start: Boolean;
              signal Xentry_296_symbol: Boolean;
              signal Xexit_297_symbol: Boolean;
              signal rr_298_symbol : Boolean;
              signal ra_299_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_295_start <= Xentry_293_symbol; -- control passed to block
              Xentry_296_symbol  <= word_access_0_295_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/$entry
              rr_298_symbol <= Xentry_296_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/rr
              ptr_deref_110_store_0_req_0 <= rr_298_symbol; -- link to DP
              ra_299_symbol <= ptr_deref_110_store_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/ra
              Xexit_297_symbol <= ra_299_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0/$exit
              word_access_0_295_symbol <= Xexit_297_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/word_access_0
            Xexit_294_symbol <= word_access_0_295_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access/$exit
            word_access_292_symbol <= Xexit_294_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/word_access
          Xexit_289_symbol <= word_access_292_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request/$exit
          ptr_deref_110_request_287_symbol <= Xexit_289_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_request
        ptr_deref_110_complete_300: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete 
          signal ptr_deref_110_complete_300_start: Boolean;
          signal Xentry_301_symbol: Boolean;
          signal Xexit_302_symbol: Boolean;
          signal word_access_303_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_110_complete_300_start <= ptr_deref_110_active_x_x266_symbol; -- control passed to block
          Xentry_301_symbol  <= ptr_deref_110_complete_300_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/$entry
          word_access_303: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access 
            signal word_access_303_start: Boolean;
            signal Xentry_304_symbol: Boolean;
            signal Xexit_305_symbol: Boolean;
            signal word_access_0_306_symbol : Boolean;
            -- 
          begin -- 
            word_access_303_start <= Xentry_301_symbol; -- control passed to block
            Xentry_304_symbol  <= word_access_303_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/$entry
            word_access_0_306: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0 
              signal word_access_0_306_start: Boolean;
              signal Xentry_307_symbol: Boolean;
              signal Xexit_308_symbol: Boolean;
              signal cr_309_symbol : Boolean;
              signal ca_310_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_306_start <= Xentry_304_symbol; -- control passed to block
              Xentry_307_symbol  <= word_access_0_306_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/$entry
              cr_309_symbol <= Xentry_307_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/cr
              ptr_deref_110_store_0_req_1 <= cr_309_symbol; -- link to DP
              ca_310_symbol <= ptr_deref_110_store_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/ca
              Xexit_308_symbol <= ca_310_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0/$exit
              word_access_0_306_symbol <= Xexit_308_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/word_access_0
            Xexit_305_symbol <= word_access_0_306_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access/$exit
            word_access_303_symbol <= Xexit_305_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/word_access
          Xexit_302_symbol <= word_access_303_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete/$exit
          ptr_deref_110_complete_300_symbol <= Xexit_302_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_110_complete
        assign_stmt_116_active_x_x311_symbol <= ptr_deref_115_complete_329_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_116_active_
        assign_stmt_116_completed_x_x312_symbol <= assign_stmt_116_active_x_x311_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_116_completed_
        ptr_deref_115_trigger_x_x313_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_trigger_ 
          signal ptr_deref_115_trigger_x_x313_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_115_trigger_x_x313_predecessors(0) <= ptr_deref_115_word_address_calculated_317_symbol;
          ptr_deref_115_trigger_x_x313_predecessors(1) <= ptr_deref_79_active_x_x62_symbol;
          ptr_deref_115_trigger_x_x313_join: join -- 
            port map( -- 
              preds => ptr_deref_115_trigger_x_x313_predecessors,
              symbol_out => ptr_deref_115_trigger_x_x313_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_trigger_
        ptr_deref_115_active_x_x314_symbol <= ptr_deref_115_request_318_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_active_
        ptr_deref_115_base_address_calculated_315_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_base_address_calculated
        ptr_deref_115_root_address_calculated_316_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_root_address_calculated
        ptr_deref_115_word_address_calculated_317_symbol <= ptr_deref_115_root_address_calculated_316_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_word_address_calculated
        ptr_deref_115_request_318: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request 
          signal ptr_deref_115_request_318_start: Boolean;
          signal Xentry_319_symbol: Boolean;
          signal Xexit_320_symbol: Boolean;
          signal word_access_321_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_115_request_318_start <= ptr_deref_115_trigger_x_x313_symbol; -- control passed to block
          Xentry_319_symbol  <= ptr_deref_115_request_318_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/$entry
          word_access_321: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access 
            signal word_access_321_start: Boolean;
            signal Xentry_322_symbol: Boolean;
            signal Xexit_323_symbol: Boolean;
            signal word_access_0_324_symbol : Boolean;
            -- 
          begin -- 
            word_access_321_start <= Xentry_319_symbol; -- control passed to block
            Xentry_322_symbol  <= word_access_321_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/$entry
            word_access_0_324: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0 
              signal word_access_0_324_start: Boolean;
              signal Xentry_325_symbol: Boolean;
              signal Xexit_326_symbol: Boolean;
              signal rr_327_symbol : Boolean;
              signal ra_328_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_324_start <= Xentry_322_symbol; -- control passed to block
              Xentry_325_symbol  <= word_access_0_324_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/$entry
              rr_327_symbol <= Xentry_325_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/rr
              ptr_deref_115_load_0_req_0 <= rr_327_symbol; -- link to DP
              ra_328_symbol <= ptr_deref_115_load_0_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/ra
              Xexit_326_symbol <= ra_328_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0/$exit
              word_access_0_324_symbol <= Xexit_326_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/word_access_0
            Xexit_323_symbol <= word_access_0_324_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access/$exit
            word_access_321_symbol <= Xexit_323_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/word_access
          Xexit_320_symbol <= word_access_321_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request/$exit
          ptr_deref_115_request_318_symbol <= Xexit_320_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_request
        ptr_deref_115_complete_329: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete 
          signal ptr_deref_115_complete_329_start: Boolean;
          signal Xentry_330_symbol: Boolean;
          signal Xexit_331_symbol: Boolean;
          signal word_access_332_symbol : Boolean;
          signal merge_req_340_symbol : Boolean;
          signal merge_ack_341_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_115_complete_329_start <= ptr_deref_115_active_x_x314_symbol; -- control passed to block
          Xentry_330_symbol  <= ptr_deref_115_complete_329_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/$entry
          word_access_332: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access 
            signal word_access_332_start: Boolean;
            signal Xentry_333_symbol: Boolean;
            signal Xexit_334_symbol: Boolean;
            signal word_access_0_335_symbol : Boolean;
            -- 
          begin -- 
            word_access_332_start <= Xentry_330_symbol; -- control passed to block
            Xentry_333_symbol  <= word_access_332_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/$entry
            word_access_0_335: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0 
              signal word_access_0_335_start: Boolean;
              signal Xentry_336_symbol: Boolean;
              signal Xexit_337_symbol: Boolean;
              signal cr_338_symbol : Boolean;
              signal ca_339_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_335_start <= Xentry_333_symbol; -- control passed to block
              Xentry_336_symbol  <= word_access_0_335_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/$entry
              cr_338_symbol <= Xentry_336_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/cr
              ptr_deref_115_load_0_req_1 <= cr_338_symbol; -- link to DP
              ca_339_symbol <= ptr_deref_115_load_0_ack_1; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/ca
              Xexit_337_symbol <= ca_339_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0/$exit
              word_access_0_335_symbol <= Xexit_337_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/word_access_0
            Xexit_334_symbol <= word_access_0_335_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access/$exit
            word_access_332_symbol <= Xexit_334_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/word_access
          merge_req_340_symbol <= word_access_332_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/merge_req
          ptr_deref_115_gather_scatter_req_0 <= merge_req_340_symbol; -- link to DP
          merge_ack_341_symbol <= ptr_deref_115_gather_scatter_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/merge_ack
          Xexit_331_symbol <= merge_ack_341_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete/$exit
          ptr_deref_115_complete_329_symbol <= Xexit_331_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/ptr_deref_115_complete
        assign_stmt_120_active_x_x342_symbol <= type_cast_119_complete_347_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_120_active_
        assign_stmt_120_completed_x_x343_symbol <= assign_stmt_120_active_x_x342_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/assign_stmt_120_completed_
        type_cast_119_active_x_x344_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_active_ 
          signal type_cast_119_active_x_x344_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_119_active_x_x344_predecessors(0) <= type_cast_119_trigger_x_x345_symbol;
          type_cast_119_active_x_x344_predecessors(1) <= simple_obj_ref_118_complete_346_symbol;
          type_cast_119_active_x_x344_join: join -- 
            port map( -- 
              preds => type_cast_119_active_x_x344_predecessors,
              symbol_out => type_cast_119_active_x_x344_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_active_
        type_cast_119_trigger_x_x345_symbol <= Xentry_46_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_trigger_
        simple_obj_ref_118_complete_346_symbol <= assign_stmt_116_completed_x_x312_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/simple_obj_ref_118_complete
        type_cast_119_complete_347: Block -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete 
          signal type_cast_119_complete_347_start: Boolean;
          signal Xentry_348_symbol: Boolean;
          signal Xexit_349_symbol: Boolean;
          signal req_350_symbol : Boolean;
          signal ack_351_symbol : Boolean;
          -- 
        begin -- 
          type_cast_119_complete_347_start <= type_cast_119_active_x_x344_symbol; -- control passed to block
          Xentry_348_symbol  <= type_cast_119_complete_347_start; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/$entry
          req_350_symbol <= Xentry_348_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/req
          type_cast_119_inst_req_0 <= req_350_symbol; -- link to DP
          ack_351_symbol <= type_cast_119_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/ack
          Xexit_349_symbol <= ack_351_symbol; -- transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete/$exit
          type_cast_119_complete_347_symbol <= Xexit_349_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/type_cast_119_complete
        Xexit_47_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/$exit 
          signal Xexit_47_predecessors: BooleanArray(6 downto 0);
          -- 
        begin -- 
          Xexit_47_predecessors(0) <= assign_stmt_81_completed_x_x59_symbol;
          Xexit_47_predecessors(1) <= ptr_deref_79_base_address_calculated_63_symbol;
          Xexit_47_predecessors(2) <= ptr_deref_84_base_address_calculated_94_symbol;
          Xexit_47_predecessors(3) <= ptr_deref_102_base_address_calculated_210_symbol;
          Xexit_47_predecessors(4) <= assign_stmt_112_completed_x_x263_symbol;
          Xexit_47_predecessors(5) <= ptr_deref_115_base_address_calculated_315_symbol;
          Xexit_47_predecessors(6) <= assign_stmt_120_completed_x_x343_symbol;
          Xexit_47_join: join -- 
            port map( -- 
              preds => Xexit_47_predecessors,
              symbol_out => Xexit_47_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125/$exit
        assign_stmt_77_to_assign_stmt_125_45_symbol <= Xexit_47_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_77_to_assign_stmt_125
      assign_stmt_129_352: Block -- branch_block_stmt_56/assign_stmt_129 
        signal assign_stmt_129_352_start: Boolean;
        signal Xentry_353_symbol: Boolean;
        signal Xexit_354_symbol: Boolean;
        signal assign_stmt_129_active_x_x355_symbol : Boolean;
        signal assign_stmt_129_completed_x_x356_symbol : Boolean;
        signal type_cast_128_active_x_x357_symbol : Boolean;
        signal type_cast_128_trigger_x_x358_symbol : Boolean;
        signal simple_obj_ref_127_complete_359_symbol : Boolean;
        signal type_cast_128_complete_360_symbol : Boolean;
        signal simple_obj_ref_126_trigger_x_x365_symbol : Boolean;
        signal simple_obj_ref_126_complete_366_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_129_352_start <= assign_stmt_129_x_xentry_x_xx_x18_symbol; -- control passed to block
        Xentry_353_symbol  <= assign_stmt_129_352_start; -- transition branch_block_stmt_56/assign_stmt_129/$entry
        assign_stmt_129_active_x_x355_symbol <= type_cast_128_complete_360_symbol; -- transition branch_block_stmt_56/assign_stmt_129/assign_stmt_129_active_
        assign_stmt_129_completed_x_x356_symbol <= simple_obj_ref_126_complete_366_symbol; -- transition branch_block_stmt_56/assign_stmt_129/assign_stmt_129_completed_
        type_cast_128_active_x_x357_block : Block -- non-trivial join transition branch_block_stmt_56/assign_stmt_129/type_cast_128_active_ 
          signal type_cast_128_active_x_x357_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_128_active_x_x357_predecessors(0) <= type_cast_128_trigger_x_x358_symbol;
          type_cast_128_active_x_x357_predecessors(1) <= simple_obj_ref_127_complete_359_symbol;
          type_cast_128_active_x_x357_join: join -- 
            port map( -- 
              preds => type_cast_128_active_x_x357_predecessors,
              symbol_out => type_cast_128_active_x_x357_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_56/assign_stmt_129/type_cast_128_active_
        type_cast_128_trigger_x_x358_symbol <= Xentry_353_symbol; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_trigger_
        simple_obj_ref_127_complete_359_symbol <= Xentry_353_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_127_complete
        type_cast_128_complete_360: Block -- branch_block_stmt_56/assign_stmt_129/type_cast_128_complete 
          signal type_cast_128_complete_360_start: Boolean;
          signal Xentry_361_symbol: Boolean;
          signal Xexit_362_symbol: Boolean;
          signal req_363_symbol : Boolean;
          signal ack_364_symbol : Boolean;
          -- 
        begin -- 
          type_cast_128_complete_360_start <= type_cast_128_active_x_x357_symbol; -- control passed to block
          Xentry_361_symbol  <= type_cast_128_complete_360_start; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/$entry
          req_363_symbol <= Xentry_361_symbol; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/req
          type_cast_128_inst_req_0 <= req_363_symbol; -- link to DP
          ack_364_symbol <= type_cast_128_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/ack
          Xexit_362_symbol <= ack_364_symbol; -- transition branch_block_stmt_56/assign_stmt_129/type_cast_128_complete/$exit
          type_cast_128_complete_360_symbol <= Xexit_362_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_129/type_cast_128_complete
        simple_obj_ref_126_trigger_x_x365_symbol <= assign_stmt_129_active_x_x355_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_trigger_
        simple_obj_ref_126_complete_366: Block -- branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete 
          signal simple_obj_ref_126_complete_366_start: Boolean;
          signal Xentry_367_symbol: Boolean;
          signal Xexit_368_symbol: Boolean;
          signal pipe_wreq_369_symbol : Boolean;
          signal pipe_wack_370_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_126_complete_366_start <= simple_obj_ref_126_trigger_x_x365_symbol; -- control passed to block
          Xentry_367_symbol  <= simple_obj_ref_126_complete_366_start; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/$entry
          pipe_wreq_369_symbol <= Xentry_367_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/pipe_wreq
          simple_obj_ref_126_inst_req_0 <= pipe_wreq_369_symbol; -- link to DP
          pipe_wack_370_symbol <= simple_obj_ref_126_inst_ack_0; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/pipe_wack
          Xexit_368_symbol <= pipe_wack_370_symbol; -- transition branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete/$exit
          simple_obj_ref_126_complete_366_symbol <= Xexit_368_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_56/assign_stmt_129/simple_obj_ref_126_complete
        Xexit_354_symbol <= assign_stmt_129_completed_x_x356_symbol; -- transition branch_block_stmt_56/assign_stmt_129/$exit
        assign_stmt_129_352_symbol <= Xexit_354_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/assign_stmt_129
      bb_0_bb_1_PhiReq_371: Block -- branch_block_stmt_56/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_371_start: Boolean;
        signal Xentry_372_symbol: Boolean;
        signal Xexit_373_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_371_start <= bb_0_bb_1_10_symbol; -- control passed to block
        Xentry_372_symbol  <= bb_0_bb_1_PhiReq_371_start; -- transition branch_block_stmt_56/bb_0_bb_1_PhiReq/$entry
        Xexit_373_symbol <= Xentry_372_symbol; -- transition branch_block_stmt_56/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_371_symbol <= Xexit_373_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/bb_0_bb_1_PhiReq
      bb_1_bb_1_PhiReq_374: Block -- branch_block_stmt_56/bb_1_bb_1_PhiReq 
        signal bb_1_bb_1_PhiReq_374_start: Boolean;
        signal Xentry_375_symbol: Boolean;
        signal Xexit_376_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_1_PhiReq_374_start <= bb_1_bb_1_20_symbol; -- control passed to block
        Xentry_375_symbol  <= bb_1_bb_1_PhiReq_374_start; -- transition branch_block_stmt_56/bb_1_bb_1_PhiReq/$entry
        Xexit_376_symbol <= Xentry_375_symbol; -- transition branch_block_stmt_56/bb_1_bb_1_PhiReq/$exit
        bb_1_bb_1_PhiReq_374_symbol <= Xexit_376_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/bb_1_bb_1_PhiReq
      merge_stmt_63_PhiReqMerge_377_symbol  <=  bb_0_bb_1_PhiReq_371_symbol or bb_1_bb_1_PhiReq_374_symbol; -- place branch_block_stmt_56/merge_stmt_63_PhiReqMerge (optimized away) 
      merge_stmt_63_PhiAck_378: Block -- branch_block_stmt_56/merge_stmt_63_PhiAck 
        signal merge_stmt_63_PhiAck_378_start: Boolean;
        signal Xentry_379_symbol: Boolean;
        signal Xexit_380_symbol: Boolean;
        signal dummy_381_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_63_PhiAck_378_start <= merge_stmt_63_PhiReqMerge_377_symbol; -- control passed to block
        Xentry_379_symbol  <= merge_stmt_63_PhiAck_378_start; -- transition branch_block_stmt_56/merge_stmt_63_PhiAck/$entry
        dummy_381_symbol <= Xentry_379_symbol; -- transition branch_block_stmt_56/merge_stmt_63_PhiAck/dummy
        Xexit_380_symbol <= dummy_381_symbol; -- transition branch_block_stmt_56/merge_stmt_63_PhiAck/$exit
        merge_stmt_63_PhiAck_378_symbol <= Xexit_380_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_56/merge_stmt_63_PhiAck
      Xexit_5_symbol <= branch_block_stmt_56_x_xexit_x_xx_x7_symbol; -- transition branch_block_stmt_56/$exit
      branch_block_stmt_56_3_symbol <= Xexit_5_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_56
    Xexit_2_symbol <= branch_block_stmt_56_3_symbol; -- transition $exit
    fin  <=  '1' when Xexit_2_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_107_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_107_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_107_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_89_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_89_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_89_root_address : std_logic_vector(2 downto 0);
    signal expr_96_wire_constant : std_logic_vector(31 downto 0);
    signal iNsTr_10_108 : std_logic_vector(31 downto 0);
    signal iNsTr_12_116 : std_logic_vector(31 downto 0);
    signal iNsTr_13_120 : std_logic_vector(31 downto 0);
    signal iNsTr_14_125 : std_logic_vector(31 downto 0);
    signal iNsTr_1_68 : std_logic_vector(31 downto 0);
    signal iNsTr_2_73 : std_logic_vector(31 downto 0);
    signal iNsTr_3_77 : std_logic_vector(31 downto 0);
    signal iNsTr_5_85 : std_logic_vector(31 downto 0);
    signal iNsTr_6_90 : std_logic_vector(31 downto 0);
    signal iNsTr_7_94 : std_logic_vector(31 downto 0);
    signal iNsTr_8_99 : std_logic_vector(31 downto 0);
    signal iNsTr_9_103 : std_logic_vector(31 downto 0);
    signal lptr_61 : std_logic_vector(31 downto 0);
    signal ptr_deref_102_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_102_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_110_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_110_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_110_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_110_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_110_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_110_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_115_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_115_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_79_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_79_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_79_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_84_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_84_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_93_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_93_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_93_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_93_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_93_word_offset_0 : std_logic_vector(2 downto 0);
    signal simple_obj_ref_71_wire : std_logic_vector(31 downto 0);
    signal type_cast_128_wire : std_logic_vector(31 downto 0);
    signal xxfooxxbodyxxlptr_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_107_final_offset <= "001";
    array_obj_ref_89_final_offset <= "001";
    expr_96_wire_constant <= "00000000000000000000000000000010";
    iNsTr_14_125 <= "00000000000000000000000000000000";
    iNsTr_1_68 <= "00000000000000000000000000000000";
    lptr_61 <= "00000000000000000000000000000000";
    ptr_deref_102_word_address_0 <= "0";
    ptr_deref_110_word_offset_0 <= "000";
    ptr_deref_115_word_address_0 <= "0";
    ptr_deref_79_word_address_0 <= "0";
    ptr_deref_84_word_address_0 <= "0";
    ptr_deref_93_word_offset_0 <= "000";
    xxfooxxbodyxxlptr_alloc_base_address <= "0";
    array_obj_ref_107_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_9_103, dout => array_obj_ref_107_resized_base_address, req => array_obj_ref_107_base_resize_req_0, ack => array_obj_ref_107_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_107_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_107_root_address, dout => iNsTr_10_108, req => array_obj_ref_107_final_reg_req_0, ack => array_obj_ref_107_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_89_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_5_85, dout => array_obj_ref_89_resized_base_address, req => array_obj_ref_89_base_resize_req_0, ack => array_obj_ref_89_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_89_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_89_root_address, dout => iNsTr_6_90, req => array_obj_ref_89_final_reg_req_0, ack => array_obj_ref_89_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_110_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_10_108, dout => ptr_deref_110_resized_base_address, req => ptr_deref_110_base_resize_req_0, ack => ptr_deref_110_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_93_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_6_90, dout => ptr_deref_93_resized_base_address, req => ptr_deref_93_base_resize_req_0, ack => ptr_deref_93_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_119_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_12_116, dout => iNsTr_13_120, req => type_cast_119_inst_req_0, ack => type_cast_119_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_128_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_13_120, dout => type_cast_128_wire, req => type_cast_128_inst_req_0, ack => type_cast_128_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_72_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_71_wire, dout => iNsTr_2_73, req => type_cast_72_inst_req_0, ack => type_cast_72_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_76_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_2_73, dout => iNsTr_3_77, req => type_cast_76_inst_req_0, ack => type_cast_76_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_102_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_102_gather_scatter_ack_0 <= ptr_deref_102_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_102_data_0;
      iNsTr_9_103 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_110_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_110_addr_0_ack_0 <= ptr_deref_110_addr_0_req_0;
      aggregated_sig <= ptr_deref_110_root_address;
      ptr_deref_110_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_110_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_110_gather_scatter_ack_0 <= ptr_deref_110_gather_scatter_req_0;
      aggregated_sig <= iNsTr_8_99;
      ptr_deref_110_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_110_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_110_root_address_inst_ack_0 <= ptr_deref_110_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_110_resized_base_address;
      ptr_deref_110_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_115_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_115_gather_scatter_ack_0 <= ptr_deref_115_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_115_data_0;
      iNsTr_12_116 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_79_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_79_gather_scatter_ack_0 <= ptr_deref_79_gather_scatter_req_0;
      aggregated_sig <= iNsTr_3_77;
      ptr_deref_79_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_84_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_84_gather_scatter_ack_0 <= ptr_deref_84_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_84_data_0;
      iNsTr_5_85 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_93_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_93_addr_0_ack_0 <= ptr_deref_93_addr_0_req_0;
      aggregated_sig <= ptr_deref_93_root_address;
      ptr_deref_93_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_93_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_93_gather_scatter_ack_0 <= ptr_deref_93_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_93_data_0;
      iNsTr_7_94 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_93_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_93_root_address_inst_ack_0 <= ptr_deref_93_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_93_resized_base_address;
      ptr_deref_93_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_107_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_107_resized_base_address;
      array_obj_ref_107_root_address <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_107_root_address_inst_req_0,
          ackL => array_obj_ref_107_root_address_inst_ack_0,
          reqR => array_obj_ref_107_root_address_inst_req_1,
          ackR => array_obj_ref_107_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_89_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_89_resized_base_address;
      array_obj_ref_89_root_address <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_89_root_address_inst_req_0,
          ackL => array_obj_ref_89_root_address_inst_ack_0,
          reqR => array_obj_ref_89_root_address_inst_req_1,
          ackR => array_obj_ref_89_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_98_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_7_94;
      iNsTr_8_99 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_98_inst_req_0,
          ackL => binary_98_inst_ack_0,
          reqR => binary_98_inst_req_1,
          ackR => binary_98_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared load operator group (0) : ptr_deref_102_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_102_load_0_req_0;
      ptr_deref_102_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_102_load_0_req_1;
      ptr_deref_102_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_102_word_address_0;
      ptr_deref_102_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(2),
          mack => memory_space_10_lr_ack(2),
          maddr => memory_space_10_lr_addr(2 downto 2),
          mtag => memory_space_10_lr_tag(2 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(2),
          mack => memory_space_10_lc_ack(2),
          mdata => memory_space_10_lc_data(95 downto 64),
          mtag => memory_space_10_lc_tag(2 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_115_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_115_load_0_req_0;
      ptr_deref_115_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_115_load_0_req_1;
      ptr_deref_115_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_115_word_address_0;
      ptr_deref_115_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(1),
          mack => memory_space_10_lr_ack(1),
          maddr => memory_space_10_lr_addr(1 downto 1),
          mtag => memory_space_10_lr_tag(1 downto 1),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(1),
          mack => memory_space_10_lc_ack(1),
          mdata => memory_space_10_lc_data(63 downto 32),
          mtag => memory_space_10_lc_tag(1 downto 1),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_84_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_84_load_0_req_0;
      ptr_deref_84_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_84_load_0_req_1;
      ptr_deref_84_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_84_word_address_0;
      ptr_deref_84_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(0),
          mack => memory_space_10_lr_ack(0),
          maddr => memory_space_10_lr_addr(0 downto 0),
          mtag => memory_space_10_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(0),
          mack => memory_space_10_lc_ack(0),
          mdata => memory_space_10_lc_data(31 downto 0),
          mtag => memory_space_10_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_93_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_93_load_0_req_0;
      ptr_deref_93_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_93_load_0_req_1;
      ptr_deref_93_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_93_word_address_0;
      ptr_deref_93_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 3,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(2 downto 0),
          mtag => memory_space_1_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared store operator group (0) : ptr_deref_110_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_110_store_0_req_0;
      ptr_deref_110_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_110_store_0_req_1;
      ptr_deref_110_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_110_word_address_0;
      data_in <= ptr_deref_110_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(2 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_79_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_79_store_0_req_0;
      ptr_deref_79_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_79_store_0_req_1;
      ptr_deref_79_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_79_word_address_0;
      data_in <= ptr_deref_79_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_10_sr_req(0),
          mack => memory_space_10_sr_ack(0),
          maddr => memory_space_10_sr_addr(0 downto 0),
          mdata => memory_space_10_sr_data(31 downto 0),
          mtag => memory_space_10_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_10_sc_req(0),
          mack => memory_space_10_sc_ack(0),
          mtag => memory_space_10_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : simple_obj_ref_71_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_71_inst_req_0;
      simple_obj_ref_71_inst_ack_0 <= ack(0);
      simple_obj_ref_71_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => foo_in_pipe_read_req(0),
          oack => foo_in_pipe_read_ack(0),
          odata => foo_in_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : simple_obj_ref_126_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_126_inst_req_0;
      simple_obj_ref_126_inst_ack_0 <= ack(0);
      data_in <= type_cast_128_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => foo_out_pipe_write_req(0),
          oack => foo_out_pipe_write_ack(0),
          odata => foo_out_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  RegisterBank_memory_space_10: register_bank -- 
    generic map(-- 
      num_loads => 3,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_10_lr_addr,
      lr_req_in => memory_space_10_lr_req,
      lr_ack_out => memory_space_10_lr_ack,
      lr_tag_in => memory_space_10_lr_tag,
      lc_req_in => memory_space_10_lc_req,
      lc_ack_out => memory_space_10_lc_ack,
      lc_data_out => memory_space_10_lc_data,
      lc_tag_out => memory_space_10_lc_tag,
      sr_addr_in => memory_space_10_sr_addr,
      sr_data_in => memory_space_10_sr_data,
      sr_req_in => memory_space_10_sr_req,
      sr_ack_out => memory_space_10_sr_ack,
      sr_tag_in => memory_space_10_sr_tag,
      sc_req_in=> memory_space_10_sc_req,
      sc_ack_out => memory_space_10_sc_ack,
      sc_tag_out => memory_space_10_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity free_queue_manager is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(1 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(1 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(1 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(1 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(1 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity free_queue_manager;
architecture Default of free_queue_manager is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_235_store_0_req_0 : boolean;
  signal simple_obj_ref_254_inst_req_0 : boolean;
  signal ptr_deref_263_load_0_req_1 : boolean;
  signal simple_obj_ref_282_load_0_ack_1 : boolean;
  signal ptr_deref_315_base_resize_req_0 : boolean;
  signal ptr_deref_315_base_resize_ack_0 : boolean;
  signal simple_obj_ref_289_load_0_ack_1 : boolean;
  signal simple_obj_ref_282_load_0_req_1 : boolean;
  signal array_obj_ref_311_final_reg_ack_0 : boolean;
  signal array_obj_ref_311_root_address_inst_req_0 : boolean;
  signal array_obj_ref_311_root_address_inst_ack_0 : boolean;
  signal ptr_deref_258_store_0_req_1 : boolean;
  signal ptr_deref_223_store_0_req_1 : boolean;
  signal if_stmt_274_branch_req_0 : boolean;
  signal ptr_deref_258_store_0_ack_0 : boolean;
  signal ptr_deref_285_store_0_ack_1 : boolean;
  signal ptr_deref_235_store_0_req_1 : boolean;
  signal ptr_deref_258_store_0_req_0 : boolean;
  signal if_stmt_274_branch_ack_0 : boolean;
  signal ptr_deref_223_store_0_ack_1 : boolean;
  signal ptr_deref_215_load_0_req_0 : boolean;
  signal simple_obj_ref_282_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_282_gather_scatter_req_0 : boolean;
  signal ptr_deref_258_gather_scatter_ack_0 : boolean;
  signal ptr_deref_258_gather_scatter_req_0 : boolean;
  signal ptr_deref_210_store_0_ack_1 : boolean;
  signal ptr_deref_223_store_0_ack_0 : boolean;
  signal ptr_deref_210_store_0_req_1 : boolean;
  signal ptr_deref_223_store_0_req_0 : boolean;
  signal binary_272_inst_ack_1 : boolean;
  signal binary_272_inst_req_1 : boolean;
  signal simple_obj_ref_282_load_0_ack_0 : boolean;
  signal if_stmt_274_branch_ack_1 : boolean;
  signal ptr_deref_235_gather_scatter_ack_0 : boolean;
  signal ptr_deref_285_store_0_req_1 : boolean;
  signal binary_272_inst_ack_0 : boolean;
  signal ptr_deref_215_gather_scatter_ack_0 : boolean;
  signal ptr_deref_223_gather_scatter_ack_0 : boolean;
  signal ptr_deref_223_gather_scatter_req_0 : boolean;
  signal ptr_deref_215_gather_scatter_req_0 : boolean;
  signal binary_272_inst_req_0 : boolean;
  signal ptr_deref_215_load_0_ack_1 : boolean;
  signal ptr_deref_210_store_0_ack_0 : boolean;
  signal ptr_deref_210_store_0_req_0 : boolean;
  signal simple_obj_ref_289_load_0_req_1 : boolean;
  signal ptr_deref_215_load_0_req_1 : boolean;
  signal simple_obj_ref_289_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_254_inst_ack_0 : boolean;
  signal ptr_deref_235_store_0_ack_0 : boolean;
  signal ptr_deref_210_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_282_load_0_req_0 : boolean;
  signal ptr_deref_210_gather_scatter_req_0 : boolean;
  signal ptr_deref_210_addr_0_ack_0 : boolean;
  signal ptr_deref_210_addr_0_req_0 : boolean;
  signal ptr_deref_215_load_0_ack_0 : boolean;
  signal ptr_deref_235_gather_scatter_req_0 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal ptr_deref_210_root_address_inst_ack_0 : boolean;
  signal ptr_deref_210_root_address_inst_req_0 : boolean;
  signal binary_220_inst_ack_1 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal binary_220_inst_req_1 : boolean;
  signal binary_220_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal simple_obj_ref_289_load_0_ack_0 : boolean;
  signal ptr_deref_210_base_resize_ack_0 : boolean;
  signal ptr_deref_285_store_0_ack_0 : boolean;
  signal ptr_deref_235_store_0_ack_1 : boolean;
  signal ptr_deref_285_store_0_req_0 : boolean;
  signal ptr_deref_210_base_resize_req_0 : boolean;
  signal array_obj_ref_311_final_reg_req_0 : boolean;
  signal if_stmt_298_branch_ack_0 : boolean;
  signal binary_296_inst_ack_1 : boolean;
  signal binary_296_inst_req_1 : boolean;
  signal binary_296_inst_req_0 : boolean;
  signal binary_296_inst_ack_0 : boolean;
  signal if_stmt_298_branch_ack_1 : boolean;
  signal type_cast_293_inst_ack_0 : boolean;
  signal type_cast_293_inst_req_0 : boolean;
  signal simple_obj_ref_243_store_0_ack_1 : boolean;
  signal ptr_deref_263_load_0_ack_0 : boolean;
  signal simple_obj_ref_243_store_0_req_1 : boolean;
  signal if_stmt_298_branch_req_0 : boolean;
  signal ptr_deref_285_gather_scatter_ack_0 : boolean;
  signal ptr_deref_263_load_0_req_0 : boolean;
  signal ptr_deref_285_gather_scatter_req_0 : boolean;
  signal ptr_deref_263_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_243_store_0_ack_0 : boolean;
  signal type_cast_255_inst_req_0 : boolean;
  signal ptr_deref_315_root_address_inst_req_0 : boolean;
  signal ptr_deref_315_root_address_inst_ack_0 : boolean;
  signal ptr_deref_315_gather_scatter_ack_0 : boolean;
  signal ptr_deref_315_load_0_req_0 : boolean;
  signal simple_obj_ref_317_store_0_req_0 : boolean;
  signal simple_obj_ref_317_store_0_ack_0 : boolean;
  signal ptr_deref_315_addr_0_req_0 : boolean;
  signal ptr_deref_315_addr_0_ack_0 : boolean;
  signal simple_obj_ref_317_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_317_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_306_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_306_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_306_load_0_ack_1 : boolean;
  signal simple_obj_ref_306_load_0_req_1 : boolean;
  signal ptr_deref_315_load_0_ack_0 : boolean;
  signal simple_obj_ref_317_store_0_req_1 : boolean;
  signal simple_obj_ref_317_store_0_ack_1 : boolean;
  signal ptr_deref_315_load_0_req_1 : boolean;
  signal ptr_deref_315_load_0_ack_1 : boolean;
  signal ptr_deref_315_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_289_gather_scatter_req_0 : boolean;
  signal ptr_deref_263_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_306_load_0_req_0 : boolean;
  signal simple_obj_ref_306_load_0_ack_0 : boolean;
  signal array_obj_ref_311_base_resize_req_0 : boolean;
  signal ptr_deref_263_load_0_ack_1 : boolean;
  signal array_obj_ref_311_base_resize_ack_0 : boolean;
  signal simple_obj_ref_289_load_0_req_0 : boolean;
  signal binary_220_inst_req_0 : boolean;
  signal ptr_deref_258_store_0_ack_1 : boolean;
  signal simple_obj_ref_243_store_0_req_0 : boolean;
  signal simple_obj_ref_243_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_243_gather_scatter_req_0 : boolean;
  signal ptr_deref_156_gather_scatter_req_0 : boolean;
  signal ptr_deref_156_gather_scatter_ack_0 : boolean;
  signal ptr_deref_156_store_0_req_0 : boolean;
  signal ptr_deref_156_store_0_ack_0 : boolean;
  signal ptr_deref_156_store_0_req_1 : boolean;
  signal ptr_deref_156_store_0_ack_1 : boolean;
  signal ptr_deref_163_load_0_req_0 : boolean;
  signal ptr_deref_163_load_0_ack_0 : boolean;
  signal ptr_deref_163_load_0_req_1 : boolean;
  signal ptr_deref_163_load_0_ack_1 : boolean;
  signal ptr_deref_163_gather_scatter_req_0 : boolean;
  signal ptr_deref_163_gather_scatter_ack_0 : boolean;
  signal type_cast_168_inst_req_0 : boolean;
  signal type_cast_168_inst_ack_0 : boolean;
  signal binary_171_inst_req_0 : boolean;
  signal binary_171_inst_ack_0 : boolean;
  signal binary_171_inst_req_1 : boolean;
  signal binary_171_inst_ack_1 : boolean;
  signal if_stmt_174_branch_req_0 : boolean;
  signal if_stmt_174_branch_ack_1 : boolean;
  signal if_stmt_174_branch_ack_0 : boolean;
  signal ptr_deref_183_load_0_req_0 : boolean;
  signal ptr_deref_183_load_0_ack_0 : boolean;
  signal ptr_deref_183_load_0_req_1 : boolean;
  signal ptr_deref_183_load_0_ack_1 : boolean;
  signal ptr_deref_183_gather_scatter_req_0 : boolean;
  signal ptr_deref_183_gather_scatter_ack_0 : boolean;
  signal binary_188_inst_req_0 : boolean;
  signal binary_188_inst_ack_0 : boolean;
  signal binary_188_inst_req_1 : boolean;
  signal binary_188_inst_ack_1 : boolean;
  signal array_obj_ref_192_index_0_resize_req_0 : boolean;
  signal array_obj_ref_192_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_192_index_0_scale_req_0 : boolean;
  signal array_obj_ref_192_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_192_index_0_scale_req_1 : boolean;
  signal array_obj_ref_192_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_192_offset_inst_req_0 : boolean;
  signal array_obj_ref_192_offset_inst_ack_0 : boolean;
  signal array_obj_ref_192_root_address_inst_req_0 : boolean;
  signal array_obj_ref_192_root_address_inst_ack_0 : boolean;
  signal addr_of_193_final_reg_req_0 : boolean;
  signal addr_of_193_final_reg_ack_0 : boolean;
  signal ptr_deref_197_load_0_req_0 : boolean;
  signal ptr_deref_197_load_0_ack_0 : boolean;
  signal ptr_deref_197_load_0_req_1 : boolean;
  signal ptr_deref_197_load_0_ack_1 : boolean;
  signal ptr_deref_197_gather_scatter_req_0 : boolean;
  signal ptr_deref_197_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_201_index_0_resize_req_0 : boolean;
  signal array_obj_ref_201_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_201_index_0_scale_req_0 : boolean;
  signal array_obj_ref_201_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_201_index_0_scale_req_1 : boolean;
  signal array_obj_ref_201_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_201_offset_inst_req_0 : boolean;
  signal array_obj_ref_201_offset_inst_ack_0 : boolean;
  signal array_obj_ref_201_root_address_inst_req_0 : boolean;
  signal array_obj_ref_201_root_address_inst_ack_0 : boolean;
  signal addr_of_202_final_reg_req_0 : boolean;
  signal addr_of_202_final_reg_ack_0 : boolean;
  signal array_obj_ref_207_base_resize_req_0 : boolean;
  signal array_obj_ref_207_base_resize_ack_0 : boolean;
  signal array_obj_ref_207_root_address_inst_req_0 : boolean;
  signal array_obj_ref_207_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_207_final_reg_req_0 : boolean;
  signal array_obj_ref_207_final_reg_ack_0 : boolean;
  signal ptr_deref_324_load_0_req_0 : boolean;
  signal ptr_deref_324_load_0_ack_0 : boolean;
  signal ptr_deref_324_load_0_req_1 : boolean;
  signal ptr_deref_324_load_0_ack_1 : boolean;
  signal ptr_deref_324_gather_scatter_req_0 : boolean;
  signal ptr_deref_324_gather_scatter_ack_0 : boolean;
  signal type_cast_328_inst_req_0 : boolean;
  signal type_cast_328_inst_ack_0 : boolean;
  signal type_cast_337_inst_req_0 : boolean;
  signal type_cast_337_inst_ack_0 : boolean;
  signal simple_obj_ref_335_inst_req_0 : boolean;
  signal simple_obj_ref_335_inst_ack_0 : boolean;
  signal ptr_deref_343_load_0_req_0 : boolean;
  signal ptr_deref_343_load_0_ack_0 : boolean;
  signal ptr_deref_343_load_0_req_1 : boolean;
  signal ptr_deref_343_load_0_ack_1 : boolean;
  signal ptr_deref_343_gather_scatter_req_0 : boolean;
  signal ptr_deref_343_gather_scatter_ack_0 : boolean;
  signal type_cast_347_inst_req_0 : boolean;
  signal type_cast_347_inst_ack_0 : boolean;
  signal binary_352_inst_req_0 : boolean;
  signal binary_352_inst_ack_0 : boolean;
  signal binary_352_inst_req_1 : boolean;
  signal binary_352_inst_ack_1 : boolean;
  signal if_stmt_354_branch_req_0 : boolean;
  signal if_stmt_354_branch_ack_1 : boolean;
  signal if_stmt_354_branch_ack_0 : boolean;
  signal simple_obj_ref_367_inst_req_0 : boolean;
  signal simple_obj_ref_367_inst_ack_0 : boolean;
  signal type_cast_368_inst_req_0 : boolean;
  signal type_cast_368_inst_ack_0 : boolean;
  signal type_cast_372_inst_req_0 : boolean;
  signal type_cast_372_inst_ack_0 : boolean;
  signal ptr_deref_375_gather_scatter_req_0 : boolean;
  signal ptr_deref_375_gather_scatter_ack_0 : boolean;
  signal ptr_deref_375_store_0_req_0 : boolean;
  signal ptr_deref_375_store_0_ack_0 : boolean;
  signal ptr_deref_375_store_0_req_1 : boolean;
  signal ptr_deref_375_store_0_ack_1 : boolean;
  signal simple_obj_ref_379_load_0_req_0 : boolean;
  signal simple_obj_ref_379_load_0_ack_0 : boolean;
  signal simple_obj_ref_379_load_0_req_1 : boolean;
  signal simple_obj_ref_379_load_0_ack_1 : boolean;
  signal simple_obj_ref_379_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_379_gather_scatter_ack_0 : boolean;
  signal ptr_deref_383_load_0_req_0 : boolean;
  signal ptr_deref_383_load_0_ack_0 : boolean;
  signal ptr_deref_383_load_0_req_1 : boolean;
  signal ptr_deref_383_load_0_ack_1 : boolean;
  signal ptr_deref_383_gather_scatter_req_0 : boolean;
  signal ptr_deref_383_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_388_base_resize_req_0 : boolean;
  signal array_obj_ref_388_base_resize_ack_0 : boolean;
  signal array_obj_ref_388_root_address_inst_req_0 : boolean;
  signal array_obj_ref_388_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_388_final_reg_req_0 : boolean;
  signal array_obj_ref_388_final_reg_ack_0 : boolean;
  signal ptr_deref_391_base_resize_req_0 : boolean;
  signal ptr_deref_391_base_resize_ack_0 : boolean;
  signal ptr_deref_391_root_address_inst_req_0 : boolean;
  signal ptr_deref_391_root_address_inst_ack_0 : boolean;
  signal ptr_deref_391_addr_0_req_0 : boolean;
  signal ptr_deref_391_addr_0_ack_0 : boolean;
  signal ptr_deref_391_gather_scatter_req_0 : boolean;
  signal ptr_deref_391_gather_scatter_ack_0 : boolean;
  signal ptr_deref_391_store_0_req_0 : boolean;
  signal ptr_deref_391_store_0_ack_0 : boolean;
  signal ptr_deref_391_store_0_req_1 : boolean;
  signal ptr_deref_391_store_0_ack_1 : boolean;
  signal ptr_deref_396_load_0_req_0 : boolean;
  signal ptr_deref_396_load_0_ack_0 : boolean;
  signal ptr_deref_396_load_0_req_1 : boolean;
  signal ptr_deref_396_load_0_ack_1 : boolean;
  signal ptr_deref_396_gather_scatter_req_0 : boolean;
  signal ptr_deref_396_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_398_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_398_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_398_store_0_req_0 : boolean;
  signal simple_obj_ref_398_store_0_ack_0 : boolean;
  signal simple_obj_ref_398_store_0_req_1 : boolean;
  signal simple_obj_ref_398_store_0_ack_1 : boolean;
  signal memory_space_11_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_11_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_11_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_11_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_11_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_11_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_11_lc_data : std_logic_vector(95 downto 0);
  signal memory_space_11_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_11_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_11_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_11_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_12_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_12_lr_tag : std_logic_vector(1 downto 0);
  signal memory_space_12_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_12_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_12_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_12_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_12_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_13_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_13_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_13_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_13_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_13_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_14_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_14_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_14_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_14_lr_tag : std_logic_vector(1 downto 0);
  signal memory_space_14_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_14_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_14_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_14_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_14_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_14_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_14_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_14_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_14_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_14_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_14_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_14_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  free_queue_manager_CP_382: Block -- control-path 
    signal free_queue_manager_CP_382_start: Boolean;
    signal Xentry_383_symbol: Boolean;
    signal Xexit_384_symbol: Boolean;
    signal branch_block_stmt_134_385_symbol : Boolean;
    -- 
  begin -- 
    free_queue_manager_CP_382_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_383_symbol  <= free_queue_manager_CP_382_start; -- transition $entry
    branch_block_stmt_134_385: Block -- branch_block_stmt_134 
      signal branch_block_stmt_134_385_start: Boolean;
      signal Xentry_386_symbol: Boolean;
      signal Xexit_387_symbol: Boolean;
      signal branch_block_stmt_134_x_xentry_x_xx_x388_symbol : Boolean;
      signal branch_block_stmt_134_x_xexit_x_xx_x389_symbol : Boolean;
      signal assign_stmt_142_to_assign_stmt_158_x_xentry_x_xx_x390_symbol : Boolean;
      signal assign_stmt_142_to_assign_stmt_158_x_xexit_x_xx_x391_symbol : Boolean;
      signal bb_0_bb_1_392_symbol : Boolean;
      signal merge_stmt_160_x_xexit_x_xx_x393_symbol : Boolean;
      signal assign_stmt_164_to_assign_stmt_173_x_xentry_x_xx_x394_symbol : Boolean;
      signal assign_stmt_164_to_assign_stmt_173_x_xexit_x_xx_x395_symbol : Boolean;
      signal if_stmt_174_x_xentry_x_xx_x396_symbol : Boolean;
      signal if_stmt_174_x_xexit_x_xx_x397_symbol : Boolean;
      signal merge_stmt_180_x_xentry_x_xx_x398_symbol : Boolean;
      signal merge_stmt_180_x_xexit_x_xx_x399_symbol : Boolean;
      signal assign_stmt_184_to_assign_stmt_225_x_xentry_x_xx_x400_symbol : Boolean;
      signal assign_stmt_184_to_assign_stmt_225_x_xexit_x_xx_x401_symbol : Boolean;
      signal bb_2_bb_1_402_symbol : Boolean;
      signal merge_stmt_227_x_xexit_x_xx_x403_symbol : Boolean;
      signal assign_stmt_233_to_assign_stmt_245_x_xentry_x_xx_x404_symbol : Boolean;
      signal assign_stmt_233_to_assign_stmt_245_x_xexit_x_xx_x405_symbol : Boolean;
      signal bb_3_bb_4_406_symbol : Boolean;
      signal merge_stmt_247_x_xexit_x_xx_x407_symbol : Boolean;
      signal assign_stmt_252_x_xentry_x_xx_x408_symbol : Boolean;
      signal assign_stmt_252_x_xexit_x_xx_x409_symbol : Boolean;
      signal assign_stmt_256_x_xentry_x_xx_x410_symbol : Boolean;
      signal assign_stmt_256_x_xexit_x_xx_x411_symbol : Boolean;
      signal assign_stmt_260_to_assign_stmt_273_x_xentry_x_xx_x412_symbol : Boolean;
      signal assign_stmt_260_to_assign_stmt_273_x_xexit_x_xx_x413_symbol : Boolean;
      signal if_stmt_274_x_xentry_x_xx_x414_symbol : Boolean;
      signal if_stmt_274_x_xexit_x_xx_x415_symbol : Boolean;
      signal merge_stmt_280_x_xentry_x_xx_x416_symbol : Boolean;
      signal merge_stmt_280_x_xexit_x_xx_x417_symbol : Boolean;
      signal assign_stmt_283_to_assign_stmt_297_x_xentry_x_xx_x418_symbol : Boolean;
      signal assign_stmt_283_to_assign_stmt_297_x_xexit_x_xx_x419_symbol : Boolean;
      signal if_stmt_298_x_xentry_x_xx_x420_symbol : Boolean;
      signal if_stmt_298_x_xexit_x_xx_x421_symbol : Boolean;
      signal merge_stmt_304_x_xentry_x_xx_x422_symbol : Boolean;
      signal merge_stmt_304_x_xexit_x_xx_x423_symbol : Boolean;
      signal assign_stmt_307_to_assign_stmt_319_x_xentry_x_xx_x424_symbol : Boolean;
      signal assign_stmt_307_to_assign_stmt_319_x_xexit_x_xx_x425_symbol : Boolean;
      signal bb_6_bb_7_426_symbol : Boolean;
      signal merge_stmt_321_x_xexit_x_xx_x427_symbol : Boolean;
      signal assign_stmt_325_to_assign_stmt_334_x_xentry_x_xx_x428_symbol : Boolean;
      signal assign_stmt_325_to_assign_stmt_334_x_xexit_x_xx_x429_symbol : Boolean;
      signal assign_stmt_338_x_xentry_x_xx_x430_symbol : Boolean;
      signal assign_stmt_338_x_xexit_x_xx_x431_symbol : Boolean;
      signal bb_7_bb_4_432_symbol : Boolean;
      signal merge_stmt_340_x_xexit_x_xx_x433_symbol : Boolean;
      signal assign_stmt_344_to_assign_stmt_353_x_xentry_x_xx_x434_symbol : Boolean;
      signal assign_stmt_344_to_assign_stmt_353_x_xexit_x_xx_x435_symbol : Boolean;
      signal if_stmt_354_x_xentry_x_xx_x436_symbol : Boolean;
      signal if_stmt_354_x_xexit_x_xx_x437_symbol : Boolean;
      signal merge_stmt_360_x_xentry_x_xx_x438_symbol : Boolean;
      signal merge_stmt_360_x_xexit_x_xx_x439_symbol : Boolean;
      signal assign_stmt_365_x_xentry_x_xx_x440_symbol : Boolean;
      signal assign_stmt_365_x_xexit_x_xx_x441_symbol : Boolean;
      signal assign_stmt_369_x_xentry_x_xx_x442_symbol : Boolean;
      signal assign_stmt_369_x_xexit_x_xx_x443_symbol : Boolean;
      signal assign_stmt_373_to_assign_stmt_400_x_xentry_x_xx_x444_symbol : Boolean;
      signal assign_stmt_373_to_assign_stmt_400_x_xexit_x_xx_x445_symbol : Boolean;
      signal bb_9_bb_4_446_symbol : Boolean;
      signal assign_stmt_142_to_assign_stmt_158_447_symbol : Boolean;
      signal assign_stmt_164_to_assign_stmt_173_481_symbol : Boolean;
      signal if_stmt_174_dead_link_534_symbol : Boolean;
      signal if_stmt_174_eval_test_538_symbol : Boolean;
      signal simple_obj_ref_175_place_542_symbol : Boolean;
      signal if_stmt_174_if_link_543_symbol : Boolean;
      signal if_stmt_174_else_link_547_symbol : Boolean;
      signal bb_1_bb_2_551_symbol : Boolean;
      signal bb_1_bb_3_552_symbol : Boolean;
      signal assign_stmt_184_to_assign_stmt_225_553_symbol : Boolean;
      signal assign_stmt_233_to_assign_stmt_245_850_symbol : Boolean;
      signal assign_stmt_252_914_symbol : Boolean;
      signal assign_stmt_256_917_symbol : Boolean;
      signal assign_stmt_260_to_assign_stmt_273_935_symbol : Boolean;
      signal if_stmt_274_dead_link_1023_symbol : Boolean;
      signal if_stmt_274_eval_test_1027_symbol : Boolean;
      signal simple_obj_ref_275_place_1031_symbol : Boolean;
      signal if_stmt_274_if_link_1032_symbol : Boolean;
      signal if_stmt_274_else_link_1036_symbol : Boolean;
      signal bb_4_bb_5_1040_symbol : Boolean;
      signal bb_4_bb_8_1041_symbol : Boolean;
      signal assign_stmt_283_to_assign_stmt_297_1042_symbol : Boolean;
      signal if_stmt_298_dead_link_1156_symbol : Boolean;
      signal if_stmt_298_eval_test_1160_symbol : Boolean;
      signal simple_obj_ref_299_place_1164_symbol : Boolean;
      signal if_stmt_298_if_link_1165_symbol : Boolean;
      signal if_stmt_298_else_link_1169_symbol : Boolean;
      signal bb_5_bb_6_1173_symbol : Boolean;
      signal bb_5_bb_7_1174_symbol : Boolean;
      signal assign_stmt_307_to_assign_stmt_319_1175_symbol : Boolean;
      signal assign_stmt_325_to_assign_stmt_334_1309_symbol : Boolean;
      signal assign_stmt_338_1353_symbol : Boolean;
      signal assign_stmt_344_to_assign_stmt_353_1372_symbol : Boolean;
      signal if_stmt_354_dead_link_1428_symbol : Boolean;
      signal if_stmt_354_eval_test_1432_symbol : Boolean;
      signal simple_obj_ref_355_place_1436_symbol : Boolean;
      signal if_stmt_354_if_link_1437_symbol : Boolean;
      signal if_stmt_354_else_link_1441_symbol : Boolean;
      signal bb_8_bb_9_1445_symbol : Boolean;
      signal bb_8_bb_4_1446_symbol : Boolean;
      signal assign_stmt_365_1447_symbol : Boolean;
      signal assign_stmt_369_1450_symbol : Boolean;
      signal assign_stmt_373_to_assign_stmt_400_1468_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_1707_symbol : Boolean;
      signal bb_2_bb_1_PhiReq_1710_symbol : Boolean;
      signal merge_stmt_160_PhiReqMerge_1713_symbol : Boolean;
      signal merge_stmt_160_PhiAck_1714_symbol : Boolean;
      signal merge_stmt_180_dead_link_1718_symbol : Boolean;
      signal bb_1_bb_2_PhiReq_1722_symbol : Boolean;
      signal merge_stmt_180_PhiReqMerge_1725_symbol : Boolean;
      signal merge_stmt_180_PhiAck_1726_symbol : Boolean;
      signal bb_1_bb_3_PhiReq_1730_symbol : Boolean;
      signal merge_stmt_227_PhiReqMerge_1733_symbol : Boolean;
      signal merge_stmt_227_PhiAck_1734_symbol : Boolean;
      signal bb_3_bb_4_PhiReq_1738_symbol : Boolean;
      signal bb_7_bb_4_PhiReq_1741_symbol : Boolean;
      signal bb_8_bb_4_PhiReq_1744_symbol : Boolean;
      signal bb_9_bb_4_PhiReq_1747_symbol : Boolean;
      signal merge_stmt_247_PhiReqMerge_1750_symbol : Boolean;
      signal merge_stmt_247_PhiAck_1751_symbol : Boolean;
      signal merge_stmt_280_dead_link_1755_symbol : Boolean;
      signal bb_4_bb_5_PhiReq_1759_symbol : Boolean;
      signal merge_stmt_280_PhiReqMerge_1762_symbol : Boolean;
      signal merge_stmt_280_PhiAck_1763_symbol : Boolean;
      signal merge_stmt_304_dead_link_1767_symbol : Boolean;
      signal bb_5_bb_6_PhiReq_1771_symbol : Boolean;
      signal merge_stmt_304_PhiReqMerge_1774_symbol : Boolean;
      signal merge_stmt_304_PhiAck_1775_symbol : Boolean;
      signal bb_5_bb_7_PhiReq_1779_symbol : Boolean;
      signal bb_6_bb_7_PhiReq_1782_symbol : Boolean;
      signal merge_stmt_321_PhiReqMerge_1785_symbol : Boolean;
      signal merge_stmt_321_PhiAck_1786_symbol : Boolean;
      signal bb_4_bb_8_PhiReq_1790_symbol : Boolean;
      signal merge_stmt_340_PhiReqMerge_1793_symbol : Boolean;
      signal merge_stmt_340_PhiAck_1794_symbol : Boolean;
      signal merge_stmt_360_dead_link_1798_symbol : Boolean;
      signal bb_8_bb_9_PhiReq_1802_symbol : Boolean;
      signal merge_stmt_360_PhiReqMerge_1805_symbol : Boolean;
      signal merge_stmt_360_PhiAck_1806_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_134_385_start <= Xentry_383_symbol; -- control passed to block
      Xentry_386_symbol  <= branch_block_stmt_134_385_start; -- transition branch_block_stmt_134/$entry
      branch_block_stmt_134_x_xentry_x_xx_x388_symbol  <=  Xentry_386_symbol; -- place branch_block_stmt_134/branch_block_stmt_134__entry__ (optimized away) 
      branch_block_stmt_134_x_xexit_x_xx_x389_symbol  <=   false ; -- place branch_block_stmt_134/branch_block_stmt_134__exit__ (optimized away) 
      assign_stmt_142_to_assign_stmt_158_x_xentry_x_xx_x390_symbol  <=  branch_block_stmt_134_x_xentry_x_xx_x388_symbol; -- place branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158__entry__ (optimized away) 
      assign_stmt_142_to_assign_stmt_158_x_xexit_x_xx_x391_symbol  <=  assign_stmt_142_to_assign_stmt_158_447_symbol; -- place branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158__exit__ (optimized away) 
      bb_0_bb_1_392_symbol  <=  assign_stmt_142_to_assign_stmt_158_x_xexit_x_xx_x391_symbol; -- place branch_block_stmt_134/bb_0_bb_1 (optimized away) 
      merge_stmt_160_x_xexit_x_xx_x393_symbol  <=  merge_stmt_160_PhiAck_1714_symbol; -- place branch_block_stmt_134/merge_stmt_160__exit__ (optimized away) 
      assign_stmt_164_to_assign_stmt_173_x_xentry_x_xx_x394_symbol  <=  merge_stmt_160_x_xexit_x_xx_x393_symbol; -- place branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173__entry__ (optimized away) 
      assign_stmt_164_to_assign_stmt_173_x_xexit_x_xx_x395_symbol  <=  assign_stmt_164_to_assign_stmt_173_481_symbol; -- place branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173__exit__ (optimized away) 
      if_stmt_174_x_xentry_x_xx_x396_symbol  <=  assign_stmt_164_to_assign_stmt_173_x_xexit_x_xx_x395_symbol; -- place branch_block_stmt_134/if_stmt_174__entry__ (optimized away) 
      if_stmt_174_x_xexit_x_xx_x397_symbol  <=  if_stmt_174_dead_link_534_symbol; -- place branch_block_stmt_134/if_stmt_174__exit__ (optimized away) 
      merge_stmt_180_x_xentry_x_xx_x398_symbol  <=  if_stmt_174_x_xexit_x_xx_x397_symbol; -- place branch_block_stmt_134/merge_stmt_180__entry__ (optimized away) 
      merge_stmt_180_x_xexit_x_xx_x399_symbol  <=  merge_stmt_180_dead_link_1718_symbol or merge_stmt_180_PhiAck_1726_symbol; -- place branch_block_stmt_134/merge_stmt_180__exit__ (optimized away) 
      assign_stmt_184_to_assign_stmt_225_x_xentry_x_xx_x400_symbol  <=  merge_stmt_180_x_xexit_x_xx_x399_symbol; -- place branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225__entry__ (optimized away) 
      assign_stmt_184_to_assign_stmt_225_x_xexit_x_xx_x401_symbol  <=  assign_stmt_184_to_assign_stmt_225_553_symbol; -- place branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225__exit__ (optimized away) 
      bb_2_bb_1_402_symbol  <=  assign_stmt_184_to_assign_stmt_225_x_xexit_x_xx_x401_symbol; -- place branch_block_stmt_134/bb_2_bb_1 (optimized away) 
      merge_stmt_227_x_xexit_x_xx_x403_symbol  <=  merge_stmt_227_PhiAck_1734_symbol; -- place branch_block_stmt_134/merge_stmt_227__exit__ (optimized away) 
      assign_stmt_233_to_assign_stmt_245_x_xentry_x_xx_x404_symbol  <=  merge_stmt_227_x_xexit_x_xx_x403_symbol; -- place branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245__entry__ (optimized away) 
      assign_stmt_233_to_assign_stmt_245_x_xexit_x_xx_x405_symbol  <=  assign_stmt_233_to_assign_stmt_245_850_symbol; -- place branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245__exit__ (optimized away) 
      bb_3_bb_4_406_symbol  <=  assign_stmt_233_to_assign_stmt_245_x_xexit_x_xx_x405_symbol; -- place branch_block_stmt_134/bb_3_bb_4 (optimized away) 
      merge_stmt_247_x_xexit_x_xx_x407_symbol  <=  merge_stmt_247_PhiAck_1751_symbol; -- place branch_block_stmt_134/merge_stmt_247__exit__ (optimized away) 
      assign_stmt_252_x_xentry_x_xx_x408_symbol  <=  merge_stmt_247_x_xexit_x_xx_x407_symbol; -- place branch_block_stmt_134/assign_stmt_252__entry__ (optimized away) 
      assign_stmt_252_x_xexit_x_xx_x409_symbol  <=  assign_stmt_252_914_symbol; -- place branch_block_stmt_134/assign_stmt_252__exit__ (optimized away) 
      assign_stmt_256_x_xentry_x_xx_x410_symbol  <=  assign_stmt_252_x_xexit_x_xx_x409_symbol; -- place branch_block_stmt_134/assign_stmt_256__entry__ (optimized away) 
      assign_stmt_256_x_xexit_x_xx_x411_symbol  <=  assign_stmt_256_917_symbol; -- place branch_block_stmt_134/assign_stmt_256__exit__ (optimized away) 
      assign_stmt_260_to_assign_stmt_273_x_xentry_x_xx_x412_symbol  <=  assign_stmt_256_x_xexit_x_xx_x411_symbol; -- place branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273__entry__ (optimized away) 
      assign_stmt_260_to_assign_stmt_273_x_xexit_x_xx_x413_symbol  <=  assign_stmt_260_to_assign_stmt_273_935_symbol; -- place branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273__exit__ (optimized away) 
      if_stmt_274_x_xentry_x_xx_x414_symbol  <=  assign_stmt_260_to_assign_stmt_273_x_xexit_x_xx_x413_symbol; -- place branch_block_stmt_134/if_stmt_274__entry__ (optimized away) 
      if_stmt_274_x_xexit_x_xx_x415_symbol  <=  if_stmt_274_dead_link_1023_symbol; -- place branch_block_stmt_134/if_stmt_274__exit__ (optimized away) 
      merge_stmt_280_x_xentry_x_xx_x416_symbol  <=  if_stmt_274_x_xexit_x_xx_x415_symbol; -- place branch_block_stmt_134/merge_stmt_280__entry__ (optimized away) 
      merge_stmt_280_x_xexit_x_xx_x417_symbol  <=  merge_stmt_280_dead_link_1755_symbol or merge_stmt_280_PhiAck_1763_symbol; -- place branch_block_stmt_134/merge_stmt_280__exit__ (optimized away) 
      assign_stmt_283_to_assign_stmt_297_x_xentry_x_xx_x418_symbol  <=  merge_stmt_280_x_xexit_x_xx_x417_symbol; -- place branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297__entry__ (optimized away) 
      assign_stmt_283_to_assign_stmt_297_x_xexit_x_xx_x419_symbol  <=  assign_stmt_283_to_assign_stmt_297_1042_symbol; -- place branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297__exit__ (optimized away) 
      if_stmt_298_x_xentry_x_xx_x420_symbol  <=  assign_stmt_283_to_assign_stmt_297_x_xexit_x_xx_x419_symbol; -- place branch_block_stmt_134/if_stmt_298__entry__ (optimized away) 
      if_stmt_298_x_xexit_x_xx_x421_symbol  <=  if_stmt_298_dead_link_1156_symbol; -- place branch_block_stmt_134/if_stmt_298__exit__ (optimized away) 
      merge_stmt_304_x_xentry_x_xx_x422_symbol  <=  if_stmt_298_x_xexit_x_xx_x421_symbol; -- place branch_block_stmt_134/merge_stmt_304__entry__ (optimized away) 
      merge_stmt_304_x_xexit_x_xx_x423_symbol  <=  merge_stmt_304_dead_link_1767_symbol or merge_stmt_304_PhiAck_1775_symbol; -- place branch_block_stmt_134/merge_stmt_304__exit__ (optimized away) 
      assign_stmt_307_to_assign_stmt_319_x_xentry_x_xx_x424_symbol  <=  merge_stmt_304_x_xexit_x_xx_x423_symbol; -- place branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319__entry__ (optimized away) 
      assign_stmt_307_to_assign_stmt_319_x_xexit_x_xx_x425_symbol  <=  assign_stmt_307_to_assign_stmt_319_1175_symbol; -- place branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319__exit__ (optimized away) 
      bb_6_bb_7_426_symbol  <=  assign_stmt_307_to_assign_stmt_319_x_xexit_x_xx_x425_symbol; -- place branch_block_stmt_134/bb_6_bb_7 (optimized away) 
      merge_stmt_321_x_xexit_x_xx_x427_symbol  <=  merge_stmt_321_PhiAck_1786_symbol; -- place branch_block_stmt_134/merge_stmt_321__exit__ (optimized away) 
      assign_stmt_325_to_assign_stmt_334_x_xentry_x_xx_x428_symbol  <=  merge_stmt_321_x_xexit_x_xx_x427_symbol; -- place branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334__entry__ (optimized away) 
      assign_stmt_325_to_assign_stmt_334_x_xexit_x_xx_x429_symbol  <=  assign_stmt_325_to_assign_stmt_334_1309_symbol; -- place branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334__exit__ (optimized away) 
      assign_stmt_338_x_xentry_x_xx_x430_symbol  <=  assign_stmt_325_to_assign_stmt_334_x_xexit_x_xx_x429_symbol; -- place branch_block_stmt_134/assign_stmt_338__entry__ (optimized away) 
      assign_stmt_338_x_xexit_x_xx_x431_symbol  <=  assign_stmt_338_1353_symbol; -- place branch_block_stmt_134/assign_stmt_338__exit__ (optimized away) 
      bb_7_bb_4_432_symbol  <=  assign_stmt_338_x_xexit_x_xx_x431_symbol; -- place branch_block_stmt_134/bb_7_bb_4 (optimized away) 
      merge_stmt_340_x_xexit_x_xx_x433_symbol  <=  merge_stmt_340_PhiAck_1794_symbol; -- place branch_block_stmt_134/merge_stmt_340__exit__ (optimized away) 
      assign_stmt_344_to_assign_stmt_353_x_xentry_x_xx_x434_symbol  <=  merge_stmt_340_x_xexit_x_xx_x433_symbol; -- place branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353__entry__ (optimized away) 
      assign_stmt_344_to_assign_stmt_353_x_xexit_x_xx_x435_symbol  <=  assign_stmt_344_to_assign_stmt_353_1372_symbol; -- place branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353__exit__ (optimized away) 
      if_stmt_354_x_xentry_x_xx_x436_symbol  <=  assign_stmt_344_to_assign_stmt_353_x_xexit_x_xx_x435_symbol; -- place branch_block_stmt_134/if_stmt_354__entry__ (optimized away) 
      if_stmt_354_x_xexit_x_xx_x437_symbol  <=  if_stmt_354_dead_link_1428_symbol; -- place branch_block_stmt_134/if_stmt_354__exit__ (optimized away) 
      merge_stmt_360_x_xentry_x_xx_x438_symbol  <=  if_stmt_354_x_xexit_x_xx_x437_symbol; -- place branch_block_stmt_134/merge_stmt_360__entry__ (optimized away) 
      merge_stmt_360_x_xexit_x_xx_x439_symbol  <=  merge_stmt_360_dead_link_1798_symbol or merge_stmt_360_PhiAck_1806_symbol; -- place branch_block_stmt_134/merge_stmt_360__exit__ (optimized away) 
      assign_stmt_365_x_xentry_x_xx_x440_symbol  <=  merge_stmt_360_x_xexit_x_xx_x439_symbol; -- place branch_block_stmt_134/assign_stmt_365__entry__ (optimized away) 
      assign_stmt_365_x_xexit_x_xx_x441_symbol  <=  assign_stmt_365_1447_symbol; -- place branch_block_stmt_134/assign_stmt_365__exit__ (optimized away) 
      assign_stmt_369_x_xentry_x_xx_x442_symbol  <=  assign_stmt_365_x_xexit_x_xx_x441_symbol; -- place branch_block_stmt_134/assign_stmt_369__entry__ (optimized away) 
      assign_stmt_369_x_xexit_x_xx_x443_symbol  <=  assign_stmt_369_1450_symbol; -- place branch_block_stmt_134/assign_stmt_369__exit__ (optimized away) 
      assign_stmt_373_to_assign_stmt_400_x_xentry_x_xx_x444_symbol  <=  assign_stmt_369_x_xexit_x_xx_x443_symbol; -- place branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400__entry__ (optimized away) 
      assign_stmt_373_to_assign_stmt_400_x_xexit_x_xx_x445_symbol  <=  assign_stmt_373_to_assign_stmt_400_1468_symbol; -- place branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400__exit__ (optimized away) 
      bb_9_bb_4_446_symbol  <=  assign_stmt_373_to_assign_stmt_400_x_xexit_x_xx_x445_symbol; -- place branch_block_stmt_134/bb_9_bb_4 (optimized away) 
      assign_stmt_142_to_assign_stmt_158_447: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158 
        signal assign_stmt_142_to_assign_stmt_158_447_start: Boolean;
        signal Xentry_448_symbol: Boolean;
        signal Xexit_449_symbol: Boolean;
        signal assign_stmt_158_active_x_x450_symbol : Boolean;
        signal assign_stmt_158_completed_x_x451_symbol : Boolean;
        signal ptr_deref_156_trigger_x_x452_symbol : Boolean;
        signal ptr_deref_156_active_x_x453_symbol : Boolean;
        signal ptr_deref_156_base_address_calculated_454_symbol : Boolean;
        signal ptr_deref_156_root_address_calculated_455_symbol : Boolean;
        signal ptr_deref_156_word_address_calculated_456_symbol : Boolean;
        signal ptr_deref_156_request_457_symbol : Boolean;
        signal ptr_deref_156_complete_470_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_142_to_assign_stmt_158_447_start <= assign_stmt_142_to_assign_stmt_158_x_xentry_x_xx_x390_symbol; -- control passed to block
        Xentry_448_symbol  <= assign_stmt_142_to_assign_stmt_158_447_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/$entry
        assign_stmt_158_active_x_x450_symbol <= Xentry_448_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/assign_stmt_158_active_
        assign_stmt_158_completed_x_x451_symbol <= ptr_deref_156_complete_470_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/assign_stmt_158_completed_
        ptr_deref_156_trigger_x_x452_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_trigger_ 
          signal ptr_deref_156_trigger_x_x452_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_156_trigger_x_x452_predecessors(0) <= ptr_deref_156_word_address_calculated_456_symbol;
          ptr_deref_156_trigger_x_x452_predecessors(1) <= assign_stmt_158_active_x_x450_symbol;
          ptr_deref_156_trigger_x_x452_join: join -- 
            port map( -- 
              preds => ptr_deref_156_trigger_x_x452_predecessors,
              symbol_out => ptr_deref_156_trigger_x_x452_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_trigger_
        ptr_deref_156_active_x_x453_symbol <= ptr_deref_156_request_457_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_active_
        ptr_deref_156_base_address_calculated_454_symbol <= Xentry_448_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_base_address_calculated
        ptr_deref_156_root_address_calculated_455_symbol <= Xentry_448_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_root_address_calculated
        ptr_deref_156_word_address_calculated_456_symbol <= ptr_deref_156_root_address_calculated_455_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_word_address_calculated
        ptr_deref_156_request_457: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request 
          signal ptr_deref_156_request_457_start: Boolean;
          signal Xentry_458_symbol: Boolean;
          signal Xexit_459_symbol: Boolean;
          signal split_req_460_symbol : Boolean;
          signal split_ack_461_symbol : Boolean;
          signal word_access_462_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_156_request_457_start <= ptr_deref_156_trigger_x_x452_symbol; -- control passed to block
          Xentry_458_symbol  <= ptr_deref_156_request_457_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/$entry
          split_req_460_symbol <= Xentry_458_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/split_req
          ptr_deref_156_gather_scatter_req_0 <= split_req_460_symbol; -- link to DP
          split_ack_461_symbol <= ptr_deref_156_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/split_ack
          word_access_462: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access 
            signal word_access_462_start: Boolean;
            signal Xentry_463_symbol: Boolean;
            signal Xexit_464_symbol: Boolean;
            signal word_access_0_465_symbol : Boolean;
            -- 
          begin -- 
            word_access_462_start <= split_ack_461_symbol; -- control passed to block
            Xentry_463_symbol  <= word_access_462_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/$entry
            word_access_0_465: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0 
              signal word_access_0_465_start: Boolean;
              signal Xentry_466_symbol: Boolean;
              signal Xexit_467_symbol: Boolean;
              signal rr_468_symbol : Boolean;
              signal ra_469_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_465_start <= Xentry_463_symbol; -- control passed to block
              Xentry_466_symbol  <= word_access_0_465_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/$entry
              rr_468_symbol <= Xentry_466_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/rr
              ptr_deref_156_store_0_req_0 <= rr_468_symbol; -- link to DP
              ra_469_symbol <= ptr_deref_156_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/ra
              Xexit_467_symbol <= ra_469_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0/$exit
              word_access_0_465_symbol <= Xexit_467_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/word_access_0
            Xexit_464_symbol <= word_access_0_465_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access/$exit
            word_access_462_symbol <= Xexit_464_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/word_access
          Xexit_459_symbol <= word_access_462_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request/$exit
          ptr_deref_156_request_457_symbol <= Xexit_459_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_request
        ptr_deref_156_complete_470: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete 
          signal ptr_deref_156_complete_470_start: Boolean;
          signal Xentry_471_symbol: Boolean;
          signal Xexit_472_symbol: Boolean;
          signal word_access_473_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_156_complete_470_start <= ptr_deref_156_active_x_x453_symbol; -- control passed to block
          Xentry_471_symbol  <= ptr_deref_156_complete_470_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/$entry
          word_access_473: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access 
            signal word_access_473_start: Boolean;
            signal Xentry_474_symbol: Boolean;
            signal Xexit_475_symbol: Boolean;
            signal word_access_0_476_symbol : Boolean;
            -- 
          begin -- 
            word_access_473_start <= Xentry_471_symbol; -- control passed to block
            Xentry_474_symbol  <= word_access_473_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/$entry
            word_access_0_476: Block -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0 
              signal word_access_0_476_start: Boolean;
              signal Xentry_477_symbol: Boolean;
              signal Xexit_478_symbol: Boolean;
              signal cr_479_symbol : Boolean;
              signal ca_480_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_476_start <= Xentry_474_symbol; -- control passed to block
              Xentry_477_symbol  <= word_access_0_476_start; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/$entry
              cr_479_symbol <= Xentry_477_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/cr
              ptr_deref_156_store_0_req_1 <= cr_479_symbol; -- link to DP
              ca_480_symbol <= ptr_deref_156_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/ca
              Xexit_478_symbol <= ca_480_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0/$exit
              word_access_0_476_symbol <= Xexit_478_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/word_access_0
            Xexit_475_symbol <= word_access_0_476_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access/$exit
            word_access_473_symbol <= Xexit_475_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/word_access
          Xexit_472_symbol <= word_access_473_symbol; -- transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete/$exit
          ptr_deref_156_complete_470_symbol <= Xexit_472_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/ptr_deref_156_complete
        Xexit_449_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/$exit 
          signal Xexit_449_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_449_predecessors(0) <= assign_stmt_158_completed_x_x451_symbol;
          Xexit_449_predecessors(1) <= ptr_deref_156_base_address_calculated_454_symbol;
          Xexit_449_join: join -- 
            port map( -- 
              preds => Xexit_449_predecessors,
              symbol_out => Xexit_449_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158/$exit
        assign_stmt_142_to_assign_stmt_158_447_symbol <= Xexit_449_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_142_to_assign_stmt_158
      assign_stmt_164_to_assign_stmt_173_481: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173 
        signal assign_stmt_164_to_assign_stmt_173_481_start: Boolean;
        signal Xentry_482_symbol: Boolean;
        signal Xexit_483_symbol: Boolean;
        signal assign_stmt_164_active_x_x484_symbol : Boolean;
        signal assign_stmt_164_completed_x_x485_symbol : Boolean;
        signal ptr_deref_163_trigger_x_x486_symbol : Boolean;
        signal ptr_deref_163_active_x_x487_symbol : Boolean;
        signal ptr_deref_163_base_address_calculated_488_symbol : Boolean;
        signal ptr_deref_163_root_address_calculated_489_symbol : Boolean;
        signal ptr_deref_163_word_address_calculated_490_symbol : Boolean;
        signal ptr_deref_163_request_491_symbol : Boolean;
        signal ptr_deref_163_complete_502_symbol : Boolean;
        signal assign_stmt_173_active_x_x515_symbol : Boolean;
        signal assign_stmt_173_completed_x_x516_symbol : Boolean;
        signal binary_171_active_x_x517_symbol : Boolean;
        signal binary_171_trigger_x_x518_symbol : Boolean;
        signal type_cast_168_active_x_x519_symbol : Boolean;
        signal type_cast_168_trigger_x_x520_symbol : Boolean;
        signal simple_obj_ref_167_complete_521_symbol : Boolean;
        signal type_cast_168_complete_522_symbol : Boolean;
        signal binary_171_complete_527_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_164_to_assign_stmt_173_481_start <= assign_stmt_164_to_assign_stmt_173_x_xentry_x_xx_x394_symbol; -- control passed to block
        Xentry_482_symbol  <= assign_stmt_164_to_assign_stmt_173_481_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/$entry
        assign_stmt_164_active_x_x484_symbol <= ptr_deref_163_complete_502_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_164_active_
        assign_stmt_164_completed_x_x485_symbol <= assign_stmt_164_active_x_x484_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_164_completed_
        ptr_deref_163_trigger_x_x486_symbol <= ptr_deref_163_word_address_calculated_490_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_trigger_
        ptr_deref_163_active_x_x487_symbol <= ptr_deref_163_request_491_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_active_
        ptr_deref_163_base_address_calculated_488_symbol <= Xentry_482_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_base_address_calculated
        ptr_deref_163_root_address_calculated_489_symbol <= Xentry_482_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_root_address_calculated
        ptr_deref_163_word_address_calculated_490_symbol <= ptr_deref_163_root_address_calculated_489_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_word_address_calculated
        ptr_deref_163_request_491: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request 
          signal ptr_deref_163_request_491_start: Boolean;
          signal Xentry_492_symbol: Boolean;
          signal Xexit_493_symbol: Boolean;
          signal word_access_494_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_163_request_491_start <= ptr_deref_163_trigger_x_x486_symbol; -- control passed to block
          Xentry_492_symbol  <= ptr_deref_163_request_491_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/$entry
          word_access_494: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access 
            signal word_access_494_start: Boolean;
            signal Xentry_495_symbol: Boolean;
            signal Xexit_496_symbol: Boolean;
            signal word_access_0_497_symbol : Boolean;
            -- 
          begin -- 
            word_access_494_start <= Xentry_492_symbol; -- control passed to block
            Xentry_495_symbol  <= word_access_494_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/$entry
            word_access_0_497: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0 
              signal word_access_0_497_start: Boolean;
              signal Xentry_498_symbol: Boolean;
              signal Xexit_499_symbol: Boolean;
              signal rr_500_symbol : Boolean;
              signal ra_501_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_497_start <= Xentry_495_symbol; -- control passed to block
              Xentry_498_symbol  <= word_access_0_497_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/$entry
              rr_500_symbol <= Xentry_498_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/rr
              ptr_deref_163_load_0_req_0 <= rr_500_symbol; -- link to DP
              ra_501_symbol <= ptr_deref_163_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/ra
              Xexit_499_symbol <= ra_501_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0/$exit
              word_access_0_497_symbol <= Xexit_499_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/word_access_0
            Xexit_496_symbol <= word_access_0_497_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access/$exit
            word_access_494_symbol <= Xexit_496_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/word_access
          Xexit_493_symbol <= word_access_494_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request/$exit
          ptr_deref_163_request_491_symbol <= Xexit_493_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_request
        ptr_deref_163_complete_502: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete 
          signal ptr_deref_163_complete_502_start: Boolean;
          signal Xentry_503_symbol: Boolean;
          signal Xexit_504_symbol: Boolean;
          signal word_access_505_symbol : Boolean;
          signal merge_req_513_symbol : Boolean;
          signal merge_ack_514_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_163_complete_502_start <= ptr_deref_163_active_x_x487_symbol; -- control passed to block
          Xentry_503_symbol  <= ptr_deref_163_complete_502_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/$entry
          word_access_505: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access 
            signal word_access_505_start: Boolean;
            signal Xentry_506_symbol: Boolean;
            signal Xexit_507_symbol: Boolean;
            signal word_access_0_508_symbol : Boolean;
            -- 
          begin -- 
            word_access_505_start <= Xentry_503_symbol; -- control passed to block
            Xentry_506_symbol  <= word_access_505_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/$entry
            word_access_0_508: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0 
              signal word_access_0_508_start: Boolean;
              signal Xentry_509_symbol: Boolean;
              signal Xexit_510_symbol: Boolean;
              signal cr_511_symbol : Boolean;
              signal ca_512_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_508_start <= Xentry_506_symbol; -- control passed to block
              Xentry_509_symbol  <= word_access_0_508_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/$entry
              cr_511_symbol <= Xentry_509_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/cr
              ptr_deref_163_load_0_req_1 <= cr_511_symbol; -- link to DP
              ca_512_symbol <= ptr_deref_163_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/ca
              Xexit_510_symbol <= ca_512_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0/$exit
              word_access_0_508_symbol <= Xexit_510_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/word_access_0
            Xexit_507_symbol <= word_access_0_508_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access/$exit
            word_access_505_symbol <= Xexit_507_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/word_access
          merge_req_513_symbol <= word_access_505_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/merge_req
          ptr_deref_163_gather_scatter_req_0 <= merge_req_513_symbol; -- link to DP
          merge_ack_514_symbol <= ptr_deref_163_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/merge_ack
          Xexit_504_symbol <= merge_ack_514_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete/$exit
          ptr_deref_163_complete_502_symbol <= Xexit_504_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/ptr_deref_163_complete
        assign_stmt_173_active_x_x515_symbol <= binary_171_complete_527_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_173_active_
        assign_stmt_173_completed_x_x516_symbol <= assign_stmt_173_active_x_x515_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/assign_stmt_173_completed_
        binary_171_active_x_x517_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_active_ 
          signal binary_171_active_x_x517_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_171_active_x_x517_predecessors(0) <= binary_171_trigger_x_x518_symbol;
          binary_171_active_x_x517_predecessors(1) <= type_cast_168_complete_522_symbol;
          binary_171_active_x_x517_join: join -- 
            port map( -- 
              preds => binary_171_active_x_x517_predecessors,
              symbol_out => binary_171_active_x_x517_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_active_
        binary_171_trigger_x_x518_symbol <= Xentry_482_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_trigger_
        type_cast_168_active_x_x519_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_active_ 
          signal type_cast_168_active_x_x519_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_168_active_x_x519_predecessors(0) <= type_cast_168_trigger_x_x520_symbol;
          type_cast_168_active_x_x519_predecessors(1) <= simple_obj_ref_167_complete_521_symbol;
          type_cast_168_active_x_x519_join: join -- 
            port map( -- 
              preds => type_cast_168_active_x_x519_predecessors,
              symbol_out => type_cast_168_active_x_x519_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_active_
        type_cast_168_trigger_x_x520_symbol <= Xentry_482_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_trigger_
        simple_obj_ref_167_complete_521_symbol <= assign_stmt_164_completed_x_x485_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/simple_obj_ref_167_complete
        type_cast_168_complete_522: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete 
          signal type_cast_168_complete_522_start: Boolean;
          signal Xentry_523_symbol: Boolean;
          signal Xexit_524_symbol: Boolean;
          signal req_525_symbol : Boolean;
          signal ack_526_symbol : Boolean;
          -- 
        begin -- 
          type_cast_168_complete_522_start <= type_cast_168_active_x_x519_symbol; -- control passed to block
          Xentry_523_symbol  <= type_cast_168_complete_522_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/$entry
          req_525_symbol <= Xentry_523_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/req
          type_cast_168_inst_req_0 <= req_525_symbol; -- link to DP
          ack_526_symbol <= type_cast_168_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/ack
          Xexit_524_symbol <= ack_526_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete/$exit
          type_cast_168_complete_522_symbol <= Xexit_524_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/type_cast_168_complete
        binary_171_complete_527: Block -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete 
          signal binary_171_complete_527_start: Boolean;
          signal Xentry_528_symbol: Boolean;
          signal Xexit_529_symbol: Boolean;
          signal rr_530_symbol : Boolean;
          signal ra_531_symbol : Boolean;
          signal cr_532_symbol : Boolean;
          signal ca_533_symbol : Boolean;
          -- 
        begin -- 
          binary_171_complete_527_start <= binary_171_active_x_x517_symbol; -- control passed to block
          Xentry_528_symbol  <= binary_171_complete_527_start; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/$entry
          rr_530_symbol <= Xentry_528_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/rr
          binary_171_inst_req_0 <= rr_530_symbol; -- link to DP
          ra_531_symbol <= binary_171_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/ra
          cr_532_symbol <= ra_531_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/cr
          binary_171_inst_req_1 <= cr_532_symbol; -- link to DP
          ca_533_symbol <= binary_171_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/ca
          Xexit_529_symbol <= ca_533_symbol; -- transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete/$exit
          binary_171_complete_527_symbol <= Xexit_529_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/binary_171_complete
        Xexit_483_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/$exit 
          signal Xexit_483_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_483_predecessors(0) <= ptr_deref_163_base_address_calculated_488_symbol;
          Xexit_483_predecessors(1) <= assign_stmt_173_completed_x_x516_symbol;
          Xexit_483_join: join -- 
            port map( -- 
              preds => Xexit_483_predecessors,
              symbol_out => Xexit_483_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173/$exit
        assign_stmt_164_to_assign_stmt_173_481_symbol <= Xexit_483_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_164_to_assign_stmt_173
      if_stmt_174_dead_link_534: Block -- branch_block_stmt_134/if_stmt_174_dead_link 
        signal if_stmt_174_dead_link_534_start: Boolean;
        signal Xentry_535_symbol: Boolean;
        signal Xexit_536_symbol: Boolean;
        signal dead_transition_537_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_dead_link_534_start <= if_stmt_174_x_xentry_x_xx_x396_symbol; -- control passed to block
        Xentry_535_symbol  <= if_stmt_174_dead_link_534_start; -- transition branch_block_stmt_134/if_stmt_174_dead_link/$entry
        dead_transition_537_symbol <= false;
        Xexit_536_symbol <= dead_transition_537_symbol; -- transition branch_block_stmt_134/if_stmt_174_dead_link/$exit
        if_stmt_174_dead_link_534_symbol <= Xexit_536_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_dead_link
      if_stmt_174_eval_test_538: Block -- branch_block_stmt_134/if_stmt_174_eval_test 
        signal if_stmt_174_eval_test_538_start: Boolean;
        signal Xentry_539_symbol: Boolean;
        signal Xexit_540_symbol: Boolean;
        signal branch_req_541_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_eval_test_538_start <= if_stmt_174_x_xentry_x_xx_x396_symbol; -- control passed to block
        Xentry_539_symbol  <= if_stmt_174_eval_test_538_start; -- transition branch_block_stmt_134/if_stmt_174_eval_test/$entry
        branch_req_541_symbol <= Xentry_539_symbol; -- transition branch_block_stmt_134/if_stmt_174_eval_test/branch_req
        if_stmt_174_branch_req_0 <= branch_req_541_symbol; -- link to DP
        Xexit_540_symbol <= branch_req_541_symbol; -- transition branch_block_stmt_134/if_stmt_174_eval_test/$exit
        if_stmt_174_eval_test_538_symbol <= Xexit_540_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_eval_test
      simple_obj_ref_175_place_542_symbol  <=  if_stmt_174_eval_test_538_symbol; -- place branch_block_stmt_134/simple_obj_ref_175_place (optimized away) 
      if_stmt_174_if_link_543: Block -- branch_block_stmt_134/if_stmt_174_if_link 
        signal if_stmt_174_if_link_543_start: Boolean;
        signal Xentry_544_symbol: Boolean;
        signal Xexit_545_symbol: Boolean;
        signal if_choice_transition_546_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_if_link_543_start <= simple_obj_ref_175_place_542_symbol; -- control passed to block
        Xentry_544_symbol  <= if_stmt_174_if_link_543_start; -- transition branch_block_stmt_134/if_stmt_174_if_link/$entry
        if_choice_transition_546_symbol <= if_stmt_174_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_174_if_link/if_choice_transition
        Xexit_545_symbol <= if_choice_transition_546_symbol; -- transition branch_block_stmt_134/if_stmt_174_if_link/$exit
        if_stmt_174_if_link_543_symbol <= Xexit_545_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_if_link
      if_stmt_174_else_link_547: Block -- branch_block_stmt_134/if_stmt_174_else_link 
        signal if_stmt_174_else_link_547_start: Boolean;
        signal Xentry_548_symbol: Boolean;
        signal Xexit_549_symbol: Boolean;
        signal else_choice_transition_550_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_174_else_link_547_start <= simple_obj_ref_175_place_542_symbol; -- control passed to block
        Xentry_548_symbol  <= if_stmt_174_else_link_547_start; -- transition branch_block_stmt_134/if_stmt_174_else_link/$entry
        else_choice_transition_550_symbol <= if_stmt_174_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_174_else_link/else_choice_transition
        Xexit_549_symbol <= else_choice_transition_550_symbol; -- transition branch_block_stmt_134/if_stmt_174_else_link/$exit
        if_stmt_174_else_link_547_symbol <= Xexit_549_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_174_else_link
      bb_1_bb_2_551_symbol  <=  if_stmt_174_if_link_543_symbol; -- place branch_block_stmt_134/bb_1_bb_2 (optimized away) 
      bb_1_bb_3_552_symbol  <=  if_stmt_174_else_link_547_symbol; -- place branch_block_stmt_134/bb_1_bb_3 (optimized away) 
      assign_stmt_184_to_assign_stmt_225_553: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225 
        signal assign_stmt_184_to_assign_stmt_225_553_start: Boolean;
        signal Xentry_554_symbol: Boolean;
        signal Xexit_555_symbol: Boolean;
        signal assign_stmt_184_active_x_x556_symbol : Boolean;
        signal assign_stmt_184_completed_x_x557_symbol : Boolean;
        signal ptr_deref_183_trigger_x_x558_symbol : Boolean;
        signal ptr_deref_183_active_x_x559_symbol : Boolean;
        signal ptr_deref_183_base_address_calculated_560_symbol : Boolean;
        signal ptr_deref_183_root_address_calculated_561_symbol : Boolean;
        signal ptr_deref_183_word_address_calculated_562_symbol : Boolean;
        signal ptr_deref_183_request_563_symbol : Boolean;
        signal ptr_deref_183_complete_574_symbol : Boolean;
        signal assign_stmt_189_active_x_x587_symbol : Boolean;
        signal assign_stmt_189_completed_x_x588_symbol : Boolean;
        signal binary_188_active_x_x589_symbol : Boolean;
        signal binary_188_trigger_x_x590_symbol : Boolean;
        signal simple_obj_ref_186_complete_591_symbol : Boolean;
        signal binary_188_complete_592_symbol : Boolean;
        signal assign_stmt_194_active_x_x599_symbol : Boolean;
        signal assign_stmt_194_completed_x_x600_symbol : Boolean;
        signal addr_of_193_active_x_x601_symbol : Boolean;
        signal addr_of_193_trigger_x_x602_symbol : Boolean;
        signal array_obj_ref_192_root_address_calculated_603_symbol : Boolean;
        signal array_obj_ref_192_indices_scaled_604_symbol : Boolean;
        signal array_obj_ref_192_offset_calculated_605_symbol : Boolean;
        signal array_obj_ref_192_index_computed_0_606_symbol : Boolean;
        signal array_obj_ref_192_index_resized_0_607_symbol : Boolean;
        signal simple_obj_ref_191_complete_608_symbol : Boolean;
        signal array_obj_ref_192_index_resize_0_609_symbol : Boolean;
        signal array_obj_ref_192_index_scale_0_614_symbol : Boolean;
        signal array_obj_ref_192_add_indices_621_symbol : Boolean;
        signal array_obj_ref_192_base_plus_offset_626_symbol : Boolean;
        signal addr_of_193_complete_631_symbol : Boolean;
        signal assign_stmt_198_active_x_x636_symbol : Boolean;
        signal assign_stmt_198_completed_x_x637_symbol : Boolean;
        signal ptr_deref_197_trigger_x_x638_symbol : Boolean;
        signal ptr_deref_197_active_x_x639_symbol : Boolean;
        signal ptr_deref_197_base_address_calculated_640_symbol : Boolean;
        signal ptr_deref_197_root_address_calculated_641_symbol : Boolean;
        signal ptr_deref_197_word_address_calculated_642_symbol : Boolean;
        signal ptr_deref_197_request_643_symbol : Boolean;
        signal ptr_deref_197_complete_654_symbol : Boolean;
        signal assign_stmt_203_active_x_x667_symbol : Boolean;
        signal assign_stmt_203_completed_x_x668_symbol : Boolean;
        signal addr_of_202_active_x_x669_symbol : Boolean;
        signal addr_of_202_trigger_x_x670_symbol : Boolean;
        signal array_obj_ref_201_root_address_calculated_671_symbol : Boolean;
        signal array_obj_ref_201_indices_scaled_672_symbol : Boolean;
        signal array_obj_ref_201_offset_calculated_673_symbol : Boolean;
        signal array_obj_ref_201_index_computed_0_674_symbol : Boolean;
        signal array_obj_ref_201_index_resized_0_675_symbol : Boolean;
        signal simple_obj_ref_200_complete_676_symbol : Boolean;
        signal array_obj_ref_201_index_resize_0_677_symbol : Boolean;
        signal array_obj_ref_201_index_scale_0_682_symbol : Boolean;
        signal array_obj_ref_201_add_indices_689_symbol : Boolean;
        signal array_obj_ref_201_base_plus_offset_694_symbol : Boolean;
        signal addr_of_202_complete_699_symbol : Boolean;
        signal assign_stmt_208_active_x_x704_symbol : Boolean;
        signal assign_stmt_208_completed_x_x705_symbol : Boolean;
        signal array_obj_ref_207_trigger_x_x706_symbol : Boolean;
        signal array_obj_ref_207_active_x_x707_symbol : Boolean;
        signal array_obj_ref_207_base_address_calculated_708_symbol : Boolean;
        signal array_obj_ref_207_root_address_calculated_709_symbol : Boolean;
        signal array_obj_ref_207_base_address_resized_710_symbol : Boolean;
        signal array_obj_ref_207_base_addr_resize_711_symbol : Boolean;
        signal array_obj_ref_207_base_plus_offset_716_symbol : Boolean;
        signal array_obj_ref_207_complete_721_symbol : Boolean;
        signal assign_stmt_212_active_x_x726_symbol : Boolean;
        signal assign_stmt_212_completed_x_x727_symbol : Boolean;
        signal simple_obj_ref_211_complete_728_symbol : Boolean;
        signal ptr_deref_210_trigger_x_x729_symbol : Boolean;
        signal ptr_deref_210_active_x_x730_symbol : Boolean;
        signal ptr_deref_210_base_address_calculated_731_symbol : Boolean;
        signal simple_obj_ref_209_complete_732_symbol : Boolean;
        signal ptr_deref_210_root_address_calculated_733_symbol : Boolean;
        signal ptr_deref_210_word_address_calculated_734_symbol : Boolean;
        signal ptr_deref_210_base_address_resized_735_symbol : Boolean;
        signal ptr_deref_210_base_addr_resize_736_symbol : Boolean;
        signal ptr_deref_210_base_plus_offset_741_symbol : Boolean;
        signal ptr_deref_210_word_addrgen_746_symbol : Boolean;
        signal ptr_deref_210_request_751_symbol : Boolean;
        signal ptr_deref_210_complete_764_symbol : Boolean;
        signal assign_stmt_216_active_x_x775_symbol : Boolean;
        signal assign_stmt_216_completed_x_x776_symbol : Boolean;
        signal ptr_deref_215_trigger_x_x777_symbol : Boolean;
        signal ptr_deref_215_active_x_x778_symbol : Boolean;
        signal ptr_deref_215_base_address_calculated_779_symbol : Boolean;
        signal ptr_deref_215_root_address_calculated_780_symbol : Boolean;
        signal ptr_deref_215_word_address_calculated_781_symbol : Boolean;
        signal ptr_deref_215_request_782_symbol : Boolean;
        signal ptr_deref_215_complete_793_symbol : Boolean;
        signal assign_stmt_221_active_x_x806_symbol : Boolean;
        signal assign_stmt_221_completed_x_x807_symbol : Boolean;
        signal binary_220_active_x_x808_symbol : Boolean;
        signal binary_220_trigger_x_x809_symbol : Boolean;
        signal simple_obj_ref_218_complete_810_symbol : Boolean;
        signal binary_220_complete_811_symbol : Boolean;
        signal assign_stmt_225_active_x_x818_symbol : Boolean;
        signal assign_stmt_225_completed_x_x819_symbol : Boolean;
        signal simple_obj_ref_224_complete_820_symbol : Boolean;
        signal ptr_deref_223_trigger_x_x821_symbol : Boolean;
        signal ptr_deref_223_active_x_x822_symbol : Boolean;
        signal ptr_deref_223_base_address_calculated_823_symbol : Boolean;
        signal ptr_deref_223_root_address_calculated_824_symbol : Boolean;
        signal ptr_deref_223_word_address_calculated_825_symbol : Boolean;
        signal ptr_deref_223_request_826_symbol : Boolean;
        signal ptr_deref_223_complete_839_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_184_to_assign_stmt_225_553_start <= assign_stmt_184_to_assign_stmt_225_x_xentry_x_xx_x400_symbol; -- control passed to block
        Xentry_554_symbol  <= assign_stmt_184_to_assign_stmt_225_553_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/$entry
        assign_stmt_184_active_x_x556_symbol <= ptr_deref_183_complete_574_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_184_active_
        assign_stmt_184_completed_x_x557_symbol <= assign_stmt_184_active_x_x556_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_184_completed_
        ptr_deref_183_trigger_x_x558_symbol <= ptr_deref_183_word_address_calculated_562_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_trigger_
        ptr_deref_183_active_x_x559_symbol <= ptr_deref_183_request_563_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_active_
        ptr_deref_183_base_address_calculated_560_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_base_address_calculated
        ptr_deref_183_root_address_calculated_561_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_root_address_calculated
        ptr_deref_183_word_address_calculated_562_symbol <= ptr_deref_183_root_address_calculated_561_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_word_address_calculated
        ptr_deref_183_request_563: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request 
          signal ptr_deref_183_request_563_start: Boolean;
          signal Xentry_564_symbol: Boolean;
          signal Xexit_565_symbol: Boolean;
          signal word_access_566_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_183_request_563_start <= ptr_deref_183_trigger_x_x558_symbol; -- control passed to block
          Xentry_564_symbol  <= ptr_deref_183_request_563_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/$entry
          word_access_566: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access 
            signal word_access_566_start: Boolean;
            signal Xentry_567_symbol: Boolean;
            signal Xexit_568_symbol: Boolean;
            signal word_access_0_569_symbol : Boolean;
            -- 
          begin -- 
            word_access_566_start <= Xentry_564_symbol; -- control passed to block
            Xentry_567_symbol  <= word_access_566_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/$entry
            word_access_0_569: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0 
              signal word_access_0_569_start: Boolean;
              signal Xentry_570_symbol: Boolean;
              signal Xexit_571_symbol: Boolean;
              signal rr_572_symbol : Boolean;
              signal ra_573_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_569_start <= Xentry_567_symbol; -- control passed to block
              Xentry_570_symbol  <= word_access_0_569_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/$entry
              rr_572_symbol <= Xentry_570_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/rr
              ptr_deref_183_load_0_req_0 <= rr_572_symbol; -- link to DP
              ra_573_symbol <= ptr_deref_183_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/ra
              Xexit_571_symbol <= ra_573_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0/$exit
              word_access_0_569_symbol <= Xexit_571_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/word_access_0
            Xexit_568_symbol <= word_access_0_569_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access/$exit
            word_access_566_symbol <= Xexit_568_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/word_access
          Xexit_565_symbol <= word_access_566_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request/$exit
          ptr_deref_183_request_563_symbol <= Xexit_565_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_request
        ptr_deref_183_complete_574: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete 
          signal ptr_deref_183_complete_574_start: Boolean;
          signal Xentry_575_symbol: Boolean;
          signal Xexit_576_symbol: Boolean;
          signal word_access_577_symbol : Boolean;
          signal merge_req_585_symbol : Boolean;
          signal merge_ack_586_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_183_complete_574_start <= ptr_deref_183_active_x_x559_symbol; -- control passed to block
          Xentry_575_symbol  <= ptr_deref_183_complete_574_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/$entry
          word_access_577: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access 
            signal word_access_577_start: Boolean;
            signal Xentry_578_symbol: Boolean;
            signal Xexit_579_symbol: Boolean;
            signal word_access_0_580_symbol : Boolean;
            -- 
          begin -- 
            word_access_577_start <= Xentry_575_symbol; -- control passed to block
            Xentry_578_symbol  <= word_access_577_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/$entry
            word_access_0_580: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0 
              signal word_access_0_580_start: Boolean;
              signal Xentry_581_symbol: Boolean;
              signal Xexit_582_symbol: Boolean;
              signal cr_583_symbol : Boolean;
              signal ca_584_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_580_start <= Xentry_578_symbol; -- control passed to block
              Xentry_581_symbol  <= word_access_0_580_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/$entry
              cr_583_symbol <= Xentry_581_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/cr
              ptr_deref_183_load_0_req_1 <= cr_583_symbol; -- link to DP
              ca_584_symbol <= ptr_deref_183_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/ca
              Xexit_582_symbol <= ca_584_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0/$exit
              word_access_0_580_symbol <= Xexit_582_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/word_access_0
            Xexit_579_symbol <= word_access_0_580_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access/$exit
            word_access_577_symbol <= Xexit_579_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/word_access
          merge_req_585_symbol <= word_access_577_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/merge_req
          ptr_deref_183_gather_scatter_req_0 <= merge_req_585_symbol; -- link to DP
          merge_ack_586_symbol <= ptr_deref_183_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/merge_ack
          Xexit_576_symbol <= merge_ack_586_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete/$exit
          ptr_deref_183_complete_574_symbol <= Xexit_576_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_183_complete
        assign_stmt_189_active_x_x587_symbol <= binary_188_complete_592_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_189_active_
        assign_stmt_189_completed_x_x588_symbol <= assign_stmt_189_active_x_x587_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_189_completed_
        binary_188_active_x_x589_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_active_ 
          signal binary_188_active_x_x589_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_188_active_x_x589_predecessors(0) <= binary_188_trigger_x_x590_symbol;
          binary_188_active_x_x589_predecessors(1) <= simple_obj_ref_186_complete_591_symbol;
          binary_188_active_x_x589_join: join -- 
            port map( -- 
              preds => binary_188_active_x_x589_predecessors,
              symbol_out => binary_188_active_x_x589_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_active_
        binary_188_trigger_x_x590_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_trigger_
        simple_obj_ref_186_complete_591_symbol <= assign_stmt_184_completed_x_x557_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_186_complete
        binary_188_complete_592: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete 
          signal binary_188_complete_592_start: Boolean;
          signal Xentry_593_symbol: Boolean;
          signal Xexit_594_symbol: Boolean;
          signal rr_595_symbol : Boolean;
          signal ra_596_symbol : Boolean;
          signal cr_597_symbol : Boolean;
          signal ca_598_symbol : Boolean;
          -- 
        begin -- 
          binary_188_complete_592_start <= binary_188_active_x_x589_symbol; -- control passed to block
          Xentry_593_symbol  <= binary_188_complete_592_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/$entry
          rr_595_symbol <= Xentry_593_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/rr
          binary_188_inst_req_0 <= rr_595_symbol; -- link to DP
          ra_596_symbol <= binary_188_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/ra
          cr_597_symbol <= ra_596_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/cr
          binary_188_inst_req_1 <= cr_597_symbol; -- link to DP
          ca_598_symbol <= binary_188_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/ca
          Xexit_594_symbol <= ca_598_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete/$exit
          binary_188_complete_592_symbol <= Xexit_594_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_188_complete
        assign_stmt_194_active_x_x599_symbol <= addr_of_193_complete_631_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_194_active_
        assign_stmt_194_completed_x_x600_symbol <= assign_stmt_194_active_x_x599_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_194_completed_
        addr_of_193_active_x_x601_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_active_ 
          signal addr_of_193_active_x_x601_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          addr_of_193_active_x_x601_predecessors(0) <= addr_of_193_trigger_x_x602_symbol;
          addr_of_193_active_x_x601_predecessors(1) <= array_obj_ref_192_root_address_calculated_603_symbol;
          addr_of_193_active_x_x601_join: join -- 
            port map( -- 
              preds => addr_of_193_active_x_x601_predecessors,
              symbol_out => addr_of_193_active_x_x601_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_active_
        addr_of_193_trigger_x_x602_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_trigger_
        array_obj_ref_192_root_address_calculated_603_symbol <= array_obj_ref_192_base_plus_offset_626_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_root_address_calculated
        array_obj_ref_192_indices_scaled_604_symbol <= array_obj_ref_192_index_scale_0_614_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_indices_scaled
        array_obj_ref_192_offset_calculated_605_symbol <= array_obj_ref_192_add_indices_621_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_offset_calculated
        array_obj_ref_192_index_computed_0_606_symbol <= simple_obj_ref_191_complete_608_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_computed_0
        array_obj_ref_192_index_resized_0_607_symbol <= array_obj_ref_192_index_resize_0_609_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resized_0
        simple_obj_ref_191_complete_608_symbol <= assign_stmt_189_completed_x_x588_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_191_complete
        array_obj_ref_192_index_resize_0_609: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0 
          signal array_obj_ref_192_index_resize_0_609_start: Boolean;
          signal Xentry_610_symbol: Boolean;
          signal Xexit_611_symbol: Boolean;
          signal index_resize_req_612_symbol : Boolean;
          signal index_resize_ack_613_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_index_resize_0_609_start <= array_obj_ref_192_index_computed_0_606_symbol; -- control passed to block
          Xentry_610_symbol  <= array_obj_ref_192_index_resize_0_609_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/$entry
          index_resize_req_612_symbol <= Xentry_610_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/index_resize_req
          array_obj_ref_192_index_0_resize_req_0 <= index_resize_req_612_symbol; -- link to DP
          index_resize_ack_613_symbol <= array_obj_ref_192_index_0_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/index_resize_ack
          Xexit_611_symbol <= index_resize_ack_613_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0/$exit
          array_obj_ref_192_index_resize_0_609_symbol <= Xexit_611_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_resize_0
        array_obj_ref_192_index_scale_0_614: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0 
          signal array_obj_ref_192_index_scale_0_614_start: Boolean;
          signal Xentry_615_symbol: Boolean;
          signal Xexit_616_symbol: Boolean;
          signal scale_rr_617_symbol : Boolean;
          signal scale_ra_618_symbol : Boolean;
          signal scale_cr_619_symbol : Boolean;
          signal scale_ca_620_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_index_scale_0_614_start <= array_obj_ref_192_index_resized_0_607_symbol; -- control passed to block
          Xentry_615_symbol  <= array_obj_ref_192_index_scale_0_614_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/$entry
          scale_rr_617_symbol <= Xentry_615_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_rr
          array_obj_ref_192_index_0_scale_req_0 <= scale_rr_617_symbol; -- link to DP
          scale_ra_618_symbol <= array_obj_ref_192_index_0_scale_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_ra
          scale_cr_619_symbol <= scale_ra_618_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_cr
          array_obj_ref_192_index_0_scale_req_1 <= scale_cr_619_symbol; -- link to DP
          scale_ca_620_symbol <= array_obj_ref_192_index_0_scale_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/scale_ca
          Xexit_616_symbol <= scale_ca_620_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0/$exit
          array_obj_ref_192_index_scale_0_614_symbol <= Xexit_616_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_index_scale_0
        array_obj_ref_192_add_indices_621: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices 
          signal array_obj_ref_192_add_indices_621_start: Boolean;
          signal Xentry_622_symbol: Boolean;
          signal Xexit_623_symbol: Boolean;
          signal final_index_req_624_symbol : Boolean;
          signal final_index_ack_625_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_add_indices_621_start <= array_obj_ref_192_indices_scaled_604_symbol; -- control passed to block
          Xentry_622_symbol  <= array_obj_ref_192_add_indices_621_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/$entry
          final_index_req_624_symbol <= Xentry_622_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/final_index_req
          array_obj_ref_192_offset_inst_req_0 <= final_index_req_624_symbol; -- link to DP
          final_index_ack_625_symbol <= array_obj_ref_192_offset_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/final_index_ack
          Xexit_623_symbol <= final_index_ack_625_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices/$exit
          array_obj_ref_192_add_indices_621_symbol <= Xexit_623_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_add_indices
        array_obj_ref_192_base_plus_offset_626: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset 
          signal array_obj_ref_192_base_plus_offset_626_start: Boolean;
          signal Xentry_627_symbol: Boolean;
          signal Xexit_628_symbol: Boolean;
          signal sum_rename_req_629_symbol : Boolean;
          signal sum_rename_ack_630_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_192_base_plus_offset_626_start <= array_obj_ref_192_offset_calculated_605_symbol; -- control passed to block
          Xentry_627_symbol  <= array_obj_ref_192_base_plus_offset_626_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/$entry
          sum_rename_req_629_symbol <= Xentry_627_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/sum_rename_req
          array_obj_ref_192_root_address_inst_req_0 <= sum_rename_req_629_symbol; -- link to DP
          sum_rename_ack_630_symbol <= array_obj_ref_192_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/sum_rename_ack
          Xexit_628_symbol <= sum_rename_ack_630_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset/$exit
          array_obj_ref_192_base_plus_offset_626_symbol <= Xexit_628_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_192_base_plus_offset
        addr_of_193_complete_631: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete 
          signal addr_of_193_complete_631_start: Boolean;
          signal Xentry_632_symbol: Boolean;
          signal Xexit_633_symbol: Boolean;
          signal final_reg_req_634_symbol : Boolean;
          signal final_reg_ack_635_symbol : Boolean;
          -- 
        begin -- 
          addr_of_193_complete_631_start <= addr_of_193_active_x_x601_symbol; -- control passed to block
          Xentry_632_symbol  <= addr_of_193_complete_631_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/$entry
          final_reg_req_634_symbol <= Xentry_632_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/final_reg_req
          addr_of_193_final_reg_req_0 <= final_reg_req_634_symbol; -- link to DP
          final_reg_ack_635_symbol <= addr_of_193_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/final_reg_ack
          Xexit_633_symbol <= final_reg_ack_635_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete/$exit
          addr_of_193_complete_631_symbol <= Xexit_633_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_193_complete
        assign_stmt_198_active_x_x636_symbol <= ptr_deref_197_complete_654_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_198_active_
        assign_stmt_198_completed_x_x637_symbol <= assign_stmt_198_active_x_x636_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_198_completed_
        ptr_deref_197_trigger_x_x638_symbol <= ptr_deref_197_word_address_calculated_642_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_trigger_
        ptr_deref_197_active_x_x639_symbol <= ptr_deref_197_request_643_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_active_
        ptr_deref_197_base_address_calculated_640_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_base_address_calculated
        ptr_deref_197_root_address_calculated_641_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_root_address_calculated
        ptr_deref_197_word_address_calculated_642_symbol <= ptr_deref_197_root_address_calculated_641_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_word_address_calculated
        ptr_deref_197_request_643: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request 
          signal ptr_deref_197_request_643_start: Boolean;
          signal Xentry_644_symbol: Boolean;
          signal Xexit_645_symbol: Boolean;
          signal word_access_646_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_197_request_643_start <= ptr_deref_197_trigger_x_x638_symbol; -- control passed to block
          Xentry_644_symbol  <= ptr_deref_197_request_643_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/$entry
          word_access_646: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access 
            signal word_access_646_start: Boolean;
            signal Xentry_647_symbol: Boolean;
            signal Xexit_648_symbol: Boolean;
            signal word_access_0_649_symbol : Boolean;
            -- 
          begin -- 
            word_access_646_start <= Xentry_644_symbol; -- control passed to block
            Xentry_647_symbol  <= word_access_646_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/$entry
            word_access_0_649: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0 
              signal word_access_0_649_start: Boolean;
              signal Xentry_650_symbol: Boolean;
              signal Xexit_651_symbol: Boolean;
              signal rr_652_symbol : Boolean;
              signal ra_653_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_649_start <= Xentry_647_symbol; -- control passed to block
              Xentry_650_symbol  <= word_access_0_649_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/$entry
              rr_652_symbol <= Xentry_650_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/rr
              ptr_deref_197_load_0_req_0 <= rr_652_symbol; -- link to DP
              ra_653_symbol <= ptr_deref_197_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/ra
              Xexit_651_symbol <= ra_653_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0/$exit
              word_access_0_649_symbol <= Xexit_651_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/word_access_0
            Xexit_648_symbol <= word_access_0_649_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access/$exit
            word_access_646_symbol <= Xexit_648_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/word_access
          Xexit_645_symbol <= word_access_646_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request/$exit
          ptr_deref_197_request_643_symbol <= Xexit_645_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_request
        ptr_deref_197_complete_654: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete 
          signal ptr_deref_197_complete_654_start: Boolean;
          signal Xentry_655_symbol: Boolean;
          signal Xexit_656_symbol: Boolean;
          signal word_access_657_symbol : Boolean;
          signal merge_req_665_symbol : Boolean;
          signal merge_ack_666_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_197_complete_654_start <= ptr_deref_197_active_x_x639_symbol; -- control passed to block
          Xentry_655_symbol  <= ptr_deref_197_complete_654_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/$entry
          word_access_657: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access 
            signal word_access_657_start: Boolean;
            signal Xentry_658_symbol: Boolean;
            signal Xexit_659_symbol: Boolean;
            signal word_access_0_660_symbol : Boolean;
            -- 
          begin -- 
            word_access_657_start <= Xentry_655_symbol; -- control passed to block
            Xentry_658_symbol  <= word_access_657_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/$entry
            word_access_0_660: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0 
              signal word_access_0_660_start: Boolean;
              signal Xentry_661_symbol: Boolean;
              signal Xexit_662_symbol: Boolean;
              signal cr_663_symbol : Boolean;
              signal ca_664_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_660_start <= Xentry_658_symbol; -- control passed to block
              Xentry_661_symbol  <= word_access_0_660_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/$entry
              cr_663_symbol <= Xentry_661_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/cr
              ptr_deref_197_load_0_req_1 <= cr_663_symbol; -- link to DP
              ca_664_symbol <= ptr_deref_197_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/ca
              Xexit_662_symbol <= ca_664_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0/$exit
              word_access_0_660_symbol <= Xexit_662_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/word_access_0
            Xexit_659_symbol <= word_access_0_660_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access/$exit
            word_access_657_symbol <= Xexit_659_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/word_access
          merge_req_665_symbol <= word_access_657_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/merge_req
          ptr_deref_197_gather_scatter_req_0 <= merge_req_665_symbol; -- link to DP
          merge_ack_666_symbol <= ptr_deref_197_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/merge_ack
          Xexit_656_symbol <= merge_ack_666_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete/$exit
          ptr_deref_197_complete_654_symbol <= Xexit_656_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_197_complete
        assign_stmt_203_active_x_x667_symbol <= addr_of_202_complete_699_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_203_active_
        assign_stmt_203_completed_x_x668_symbol <= assign_stmt_203_active_x_x667_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_203_completed_
        addr_of_202_active_x_x669_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_active_ 
          signal addr_of_202_active_x_x669_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          addr_of_202_active_x_x669_predecessors(0) <= addr_of_202_trigger_x_x670_symbol;
          addr_of_202_active_x_x669_predecessors(1) <= array_obj_ref_201_root_address_calculated_671_symbol;
          addr_of_202_active_x_x669_join: join -- 
            port map( -- 
              preds => addr_of_202_active_x_x669_predecessors,
              symbol_out => addr_of_202_active_x_x669_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_active_
        addr_of_202_trigger_x_x670_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_trigger_
        array_obj_ref_201_root_address_calculated_671_symbol <= array_obj_ref_201_base_plus_offset_694_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_root_address_calculated
        array_obj_ref_201_indices_scaled_672_symbol <= array_obj_ref_201_index_scale_0_682_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_indices_scaled
        array_obj_ref_201_offset_calculated_673_symbol <= array_obj_ref_201_add_indices_689_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_offset_calculated
        array_obj_ref_201_index_computed_0_674_symbol <= simple_obj_ref_200_complete_676_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_computed_0
        array_obj_ref_201_index_resized_0_675_symbol <= array_obj_ref_201_index_resize_0_677_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resized_0
        simple_obj_ref_200_complete_676_symbol <= assign_stmt_198_completed_x_x637_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_200_complete
        array_obj_ref_201_index_resize_0_677: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0 
          signal array_obj_ref_201_index_resize_0_677_start: Boolean;
          signal Xentry_678_symbol: Boolean;
          signal Xexit_679_symbol: Boolean;
          signal index_resize_req_680_symbol : Boolean;
          signal index_resize_ack_681_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_index_resize_0_677_start <= array_obj_ref_201_index_computed_0_674_symbol; -- control passed to block
          Xentry_678_symbol  <= array_obj_ref_201_index_resize_0_677_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/$entry
          index_resize_req_680_symbol <= Xentry_678_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/index_resize_req
          array_obj_ref_201_index_0_resize_req_0 <= index_resize_req_680_symbol; -- link to DP
          index_resize_ack_681_symbol <= array_obj_ref_201_index_0_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/index_resize_ack
          Xexit_679_symbol <= index_resize_ack_681_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0/$exit
          array_obj_ref_201_index_resize_0_677_symbol <= Xexit_679_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_resize_0
        array_obj_ref_201_index_scale_0_682: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0 
          signal array_obj_ref_201_index_scale_0_682_start: Boolean;
          signal Xentry_683_symbol: Boolean;
          signal Xexit_684_symbol: Boolean;
          signal scale_rr_685_symbol : Boolean;
          signal scale_ra_686_symbol : Boolean;
          signal scale_cr_687_symbol : Boolean;
          signal scale_ca_688_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_index_scale_0_682_start <= array_obj_ref_201_index_resized_0_675_symbol; -- control passed to block
          Xentry_683_symbol  <= array_obj_ref_201_index_scale_0_682_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/$entry
          scale_rr_685_symbol <= Xentry_683_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_rr
          array_obj_ref_201_index_0_scale_req_0 <= scale_rr_685_symbol; -- link to DP
          scale_ra_686_symbol <= array_obj_ref_201_index_0_scale_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_ra
          scale_cr_687_symbol <= scale_ra_686_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_cr
          array_obj_ref_201_index_0_scale_req_1 <= scale_cr_687_symbol; -- link to DP
          scale_ca_688_symbol <= array_obj_ref_201_index_0_scale_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/scale_ca
          Xexit_684_symbol <= scale_ca_688_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0/$exit
          array_obj_ref_201_index_scale_0_682_symbol <= Xexit_684_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_index_scale_0
        array_obj_ref_201_add_indices_689: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices 
          signal array_obj_ref_201_add_indices_689_start: Boolean;
          signal Xentry_690_symbol: Boolean;
          signal Xexit_691_symbol: Boolean;
          signal final_index_req_692_symbol : Boolean;
          signal final_index_ack_693_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_add_indices_689_start <= array_obj_ref_201_indices_scaled_672_symbol; -- control passed to block
          Xentry_690_symbol  <= array_obj_ref_201_add_indices_689_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/$entry
          final_index_req_692_symbol <= Xentry_690_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/final_index_req
          array_obj_ref_201_offset_inst_req_0 <= final_index_req_692_symbol; -- link to DP
          final_index_ack_693_symbol <= array_obj_ref_201_offset_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/final_index_ack
          Xexit_691_symbol <= final_index_ack_693_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices/$exit
          array_obj_ref_201_add_indices_689_symbol <= Xexit_691_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_add_indices
        array_obj_ref_201_base_plus_offset_694: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset 
          signal array_obj_ref_201_base_plus_offset_694_start: Boolean;
          signal Xentry_695_symbol: Boolean;
          signal Xexit_696_symbol: Boolean;
          signal sum_rename_req_697_symbol : Boolean;
          signal sum_rename_ack_698_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_201_base_plus_offset_694_start <= array_obj_ref_201_offset_calculated_673_symbol; -- control passed to block
          Xentry_695_symbol  <= array_obj_ref_201_base_plus_offset_694_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/$entry
          sum_rename_req_697_symbol <= Xentry_695_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/sum_rename_req
          array_obj_ref_201_root_address_inst_req_0 <= sum_rename_req_697_symbol; -- link to DP
          sum_rename_ack_698_symbol <= array_obj_ref_201_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/sum_rename_ack
          Xexit_696_symbol <= sum_rename_ack_698_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset/$exit
          array_obj_ref_201_base_plus_offset_694_symbol <= Xexit_696_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_201_base_plus_offset
        addr_of_202_complete_699: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete 
          signal addr_of_202_complete_699_start: Boolean;
          signal Xentry_700_symbol: Boolean;
          signal Xexit_701_symbol: Boolean;
          signal final_reg_req_702_symbol : Boolean;
          signal final_reg_ack_703_symbol : Boolean;
          -- 
        begin -- 
          addr_of_202_complete_699_start <= addr_of_202_active_x_x669_symbol; -- control passed to block
          Xentry_700_symbol  <= addr_of_202_complete_699_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/$entry
          final_reg_req_702_symbol <= Xentry_700_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/final_reg_req
          addr_of_202_final_reg_req_0 <= final_reg_req_702_symbol; -- link to DP
          final_reg_ack_703_symbol <= addr_of_202_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/final_reg_ack
          Xexit_701_symbol <= final_reg_ack_703_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete/$exit
          addr_of_202_complete_699_symbol <= Xexit_701_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/addr_of_202_complete
        assign_stmt_208_active_x_x704_symbol <= array_obj_ref_207_complete_721_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_208_active_
        assign_stmt_208_completed_x_x705_symbol <= assign_stmt_208_active_x_x704_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_208_completed_
        array_obj_ref_207_trigger_x_x706_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_trigger_
        array_obj_ref_207_active_x_x707_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_active_ 
          signal array_obj_ref_207_active_x_x707_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_207_active_x_x707_predecessors(0) <= array_obj_ref_207_trigger_x_x706_symbol;
          array_obj_ref_207_active_x_x707_predecessors(1) <= array_obj_ref_207_root_address_calculated_709_symbol;
          array_obj_ref_207_active_x_x707_join: join -- 
            port map( -- 
              preds => array_obj_ref_207_active_x_x707_predecessors,
              symbol_out => array_obj_ref_207_active_x_x707_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_active_
        array_obj_ref_207_base_address_calculated_708_symbol <= assign_stmt_203_completed_x_x668_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_address_calculated
        array_obj_ref_207_root_address_calculated_709_symbol <= array_obj_ref_207_base_plus_offset_716_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_root_address_calculated
        array_obj_ref_207_base_address_resized_710_symbol <= array_obj_ref_207_base_addr_resize_711_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_address_resized
        array_obj_ref_207_base_addr_resize_711: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize 
          signal array_obj_ref_207_base_addr_resize_711_start: Boolean;
          signal Xentry_712_symbol: Boolean;
          signal Xexit_713_symbol: Boolean;
          signal base_resize_req_714_symbol : Boolean;
          signal base_resize_ack_715_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_207_base_addr_resize_711_start <= array_obj_ref_207_base_address_calculated_708_symbol; -- control passed to block
          Xentry_712_symbol  <= array_obj_ref_207_base_addr_resize_711_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/$entry
          base_resize_req_714_symbol <= Xentry_712_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/base_resize_req
          array_obj_ref_207_base_resize_req_0 <= base_resize_req_714_symbol; -- link to DP
          base_resize_ack_715_symbol <= array_obj_ref_207_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/base_resize_ack
          Xexit_713_symbol <= base_resize_ack_715_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize/$exit
          array_obj_ref_207_base_addr_resize_711_symbol <= Xexit_713_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_addr_resize
        array_obj_ref_207_base_plus_offset_716: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset 
          signal array_obj_ref_207_base_plus_offset_716_start: Boolean;
          signal Xentry_717_symbol: Boolean;
          signal Xexit_718_symbol: Boolean;
          signal sum_rename_req_719_symbol : Boolean;
          signal sum_rename_ack_720_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_207_base_plus_offset_716_start <= array_obj_ref_207_base_address_resized_710_symbol; -- control passed to block
          Xentry_717_symbol  <= array_obj_ref_207_base_plus_offset_716_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/$entry
          sum_rename_req_719_symbol <= Xentry_717_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/sum_rename_req
          array_obj_ref_207_root_address_inst_req_0 <= sum_rename_req_719_symbol; -- link to DP
          sum_rename_ack_720_symbol <= array_obj_ref_207_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/sum_rename_ack
          Xexit_718_symbol <= sum_rename_ack_720_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset/$exit
          array_obj_ref_207_base_plus_offset_716_symbol <= Xexit_718_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_base_plus_offset
        array_obj_ref_207_complete_721: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete 
          signal array_obj_ref_207_complete_721_start: Boolean;
          signal Xentry_722_symbol: Boolean;
          signal Xexit_723_symbol: Boolean;
          signal final_reg_req_724_symbol : Boolean;
          signal final_reg_ack_725_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_207_complete_721_start <= array_obj_ref_207_active_x_x707_symbol; -- control passed to block
          Xentry_722_symbol  <= array_obj_ref_207_complete_721_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/$entry
          final_reg_req_724_symbol <= Xentry_722_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/final_reg_req
          array_obj_ref_207_final_reg_req_0 <= final_reg_req_724_symbol; -- link to DP
          final_reg_ack_725_symbol <= array_obj_ref_207_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/final_reg_ack
          Xexit_723_symbol <= final_reg_ack_725_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete/$exit
          array_obj_ref_207_complete_721_symbol <= Xexit_723_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/array_obj_ref_207_complete
        assign_stmt_212_active_x_x726_symbol <= simple_obj_ref_211_complete_728_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_212_active_
        assign_stmt_212_completed_x_x727_symbol <= ptr_deref_210_complete_764_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_212_completed_
        simple_obj_ref_211_complete_728_symbol <= assign_stmt_194_completed_x_x600_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_211_complete
        ptr_deref_210_trigger_x_x729_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_trigger_ 
          signal ptr_deref_210_trigger_x_x729_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          ptr_deref_210_trigger_x_x729_predecessors(0) <= ptr_deref_210_word_address_calculated_734_symbol;
          ptr_deref_210_trigger_x_x729_predecessors(1) <= ptr_deref_210_base_address_calculated_731_symbol;
          ptr_deref_210_trigger_x_x729_predecessors(2) <= assign_stmt_212_active_x_x726_symbol;
          ptr_deref_210_trigger_x_x729_join: join -- 
            port map( -- 
              preds => ptr_deref_210_trigger_x_x729_predecessors,
              symbol_out => ptr_deref_210_trigger_x_x729_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_trigger_
        ptr_deref_210_active_x_x730_symbol <= ptr_deref_210_request_751_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_active_
        ptr_deref_210_base_address_calculated_731_symbol <= simple_obj_ref_209_complete_732_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_address_calculated
        simple_obj_ref_209_complete_732_symbol <= assign_stmt_208_completed_x_x705_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_209_complete
        ptr_deref_210_root_address_calculated_733_symbol <= ptr_deref_210_base_plus_offset_741_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_root_address_calculated
        ptr_deref_210_word_address_calculated_734_symbol <= ptr_deref_210_word_addrgen_746_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_address_calculated
        ptr_deref_210_base_address_resized_735_symbol <= ptr_deref_210_base_addr_resize_736_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_address_resized
        ptr_deref_210_base_addr_resize_736: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize 
          signal ptr_deref_210_base_addr_resize_736_start: Boolean;
          signal Xentry_737_symbol: Boolean;
          signal Xexit_738_symbol: Boolean;
          signal base_resize_req_739_symbol : Boolean;
          signal base_resize_ack_740_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_base_addr_resize_736_start <= ptr_deref_210_base_address_calculated_731_symbol; -- control passed to block
          Xentry_737_symbol  <= ptr_deref_210_base_addr_resize_736_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/$entry
          base_resize_req_739_symbol <= Xentry_737_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/base_resize_req
          ptr_deref_210_base_resize_req_0 <= base_resize_req_739_symbol; -- link to DP
          base_resize_ack_740_symbol <= ptr_deref_210_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/base_resize_ack
          Xexit_738_symbol <= base_resize_ack_740_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize/$exit
          ptr_deref_210_base_addr_resize_736_symbol <= Xexit_738_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_addr_resize
        ptr_deref_210_base_plus_offset_741: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset 
          signal ptr_deref_210_base_plus_offset_741_start: Boolean;
          signal Xentry_742_symbol: Boolean;
          signal Xexit_743_symbol: Boolean;
          signal sum_rename_req_744_symbol : Boolean;
          signal sum_rename_ack_745_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_base_plus_offset_741_start <= ptr_deref_210_base_address_resized_735_symbol; -- control passed to block
          Xentry_742_symbol  <= ptr_deref_210_base_plus_offset_741_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/$entry
          sum_rename_req_744_symbol <= Xentry_742_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/sum_rename_req
          ptr_deref_210_root_address_inst_req_0 <= sum_rename_req_744_symbol; -- link to DP
          sum_rename_ack_745_symbol <= ptr_deref_210_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/sum_rename_ack
          Xexit_743_symbol <= sum_rename_ack_745_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset/$exit
          ptr_deref_210_base_plus_offset_741_symbol <= Xexit_743_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_base_plus_offset
        ptr_deref_210_word_addrgen_746: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen 
          signal ptr_deref_210_word_addrgen_746_start: Boolean;
          signal Xentry_747_symbol: Boolean;
          signal Xexit_748_symbol: Boolean;
          signal root_rename_req_749_symbol : Boolean;
          signal root_rename_ack_750_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_word_addrgen_746_start <= ptr_deref_210_root_address_calculated_733_symbol; -- control passed to block
          Xentry_747_symbol  <= ptr_deref_210_word_addrgen_746_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/$entry
          root_rename_req_749_symbol <= Xentry_747_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/root_rename_req
          ptr_deref_210_addr_0_req_0 <= root_rename_req_749_symbol; -- link to DP
          root_rename_ack_750_symbol <= ptr_deref_210_addr_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/root_rename_ack
          Xexit_748_symbol <= root_rename_ack_750_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen/$exit
          ptr_deref_210_word_addrgen_746_symbol <= Xexit_748_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_word_addrgen
        ptr_deref_210_request_751: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request 
          signal ptr_deref_210_request_751_start: Boolean;
          signal Xentry_752_symbol: Boolean;
          signal Xexit_753_symbol: Boolean;
          signal split_req_754_symbol : Boolean;
          signal split_ack_755_symbol : Boolean;
          signal word_access_756_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_request_751_start <= ptr_deref_210_trigger_x_x729_symbol; -- control passed to block
          Xentry_752_symbol  <= ptr_deref_210_request_751_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/$entry
          split_req_754_symbol <= Xentry_752_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/split_req
          ptr_deref_210_gather_scatter_req_0 <= split_req_754_symbol; -- link to DP
          split_ack_755_symbol <= ptr_deref_210_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/split_ack
          word_access_756: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access 
            signal word_access_756_start: Boolean;
            signal Xentry_757_symbol: Boolean;
            signal Xexit_758_symbol: Boolean;
            signal word_access_0_759_symbol : Boolean;
            -- 
          begin -- 
            word_access_756_start <= split_ack_755_symbol; -- control passed to block
            Xentry_757_symbol  <= word_access_756_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/$entry
            word_access_0_759: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0 
              signal word_access_0_759_start: Boolean;
              signal Xentry_760_symbol: Boolean;
              signal Xexit_761_symbol: Boolean;
              signal rr_762_symbol : Boolean;
              signal ra_763_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_759_start <= Xentry_757_symbol; -- control passed to block
              Xentry_760_symbol  <= word_access_0_759_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/$entry
              rr_762_symbol <= Xentry_760_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/rr
              ptr_deref_210_store_0_req_0 <= rr_762_symbol; -- link to DP
              ra_763_symbol <= ptr_deref_210_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/ra
              Xexit_761_symbol <= ra_763_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0/$exit
              word_access_0_759_symbol <= Xexit_761_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/word_access_0
            Xexit_758_symbol <= word_access_0_759_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access/$exit
            word_access_756_symbol <= Xexit_758_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/word_access
          Xexit_753_symbol <= word_access_756_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request/$exit
          ptr_deref_210_request_751_symbol <= Xexit_753_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_request
        ptr_deref_210_complete_764: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete 
          signal ptr_deref_210_complete_764_start: Boolean;
          signal Xentry_765_symbol: Boolean;
          signal Xexit_766_symbol: Boolean;
          signal word_access_767_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_210_complete_764_start <= ptr_deref_210_active_x_x730_symbol; -- control passed to block
          Xentry_765_symbol  <= ptr_deref_210_complete_764_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/$entry
          word_access_767: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access 
            signal word_access_767_start: Boolean;
            signal Xentry_768_symbol: Boolean;
            signal Xexit_769_symbol: Boolean;
            signal word_access_0_770_symbol : Boolean;
            -- 
          begin -- 
            word_access_767_start <= Xentry_765_symbol; -- control passed to block
            Xentry_768_symbol  <= word_access_767_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/$entry
            word_access_0_770: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0 
              signal word_access_0_770_start: Boolean;
              signal Xentry_771_symbol: Boolean;
              signal Xexit_772_symbol: Boolean;
              signal cr_773_symbol : Boolean;
              signal ca_774_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_770_start <= Xentry_768_symbol; -- control passed to block
              Xentry_771_symbol  <= word_access_0_770_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/$entry
              cr_773_symbol <= Xentry_771_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/cr
              ptr_deref_210_store_0_req_1 <= cr_773_symbol; -- link to DP
              ca_774_symbol <= ptr_deref_210_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/ca
              Xexit_772_symbol <= ca_774_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0/$exit
              word_access_0_770_symbol <= Xexit_772_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/word_access_0
            Xexit_769_symbol <= word_access_0_770_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access/$exit
            word_access_767_symbol <= Xexit_769_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/word_access
          Xexit_766_symbol <= word_access_767_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete/$exit
          ptr_deref_210_complete_764_symbol <= Xexit_766_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_210_complete
        assign_stmt_216_active_x_x775_symbol <= ptr_deref_215_complete_793_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_216_active_
        assign_stmt_216_completed_x_x776_symbol <= assign_stmt_216_active_x_x775_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_216_completed_
        ptr_deref_215_trigger_x_x777_symbol <= ptr_deref_215_word_address_calculated_781_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_trigger_
        ptr_deref_215_active_x_x778_symbol <= ptr_deref_215_request_782_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_active_
        ptr_deref_215_base_address_calculated_779_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_base_address_calculated
        ptr_deref_215_root_address_calculated_780_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_root_address_calculated
        ptr_deref_215_word_address_calculated_781_symbol <= ptr_deref_215_root_address_calculated_780_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_word_address_calculated
        ptr_deref_215_request_782: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request 
          signal ptr_deref_215_request_782_start: Boolean;
          signal Xentry_783_symbol: Boolean;
          signal Xexit_784_symbol: Boolean;
          signal word_access_785_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_215_request_782_start <= ptr_deref_215_trigger_x_x777_symbol; -- control passed to block
          Xentry_783_symbol  <= ptr_deref_215_request_782_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/$entry
          word_access_785: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access 
            signal word_access_785_start: Boolean;
            signal Xentry_786_symbol: Boolean;
            signal Xexit_787_symbol: Boolean;
            signal word_access_0_788_symbol : Boolean;
            -- 
          begin -- 
            word_access_785_start <= Xentry_783_symbol; -- control passed to block
            Xentry_786_symbol  <= word_access_785_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/$entry
            word_access_0_788: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0 
              signal word_access_0_788_start: Boolean;
              signal Xentry_789_symbol: Boolean;
              signal Xexit_790_symbol: Boolean;
              signal rr_791_symbol : Boolean;
              signal ra_792_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_788_start <= Xentry_786_symbol; -- control passed to block
              Xentry_789_symbol  <= word_access_0_788_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/$entry
              rr_791_symbol <= Xentry_789_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/rr
              ptr_deref_215_load_0_req_0 <= rr_791_symbol; -- link to DP
              ra_792_symbol <= ptr_deref_215_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/ra
              Xexit_790_symbol <= ra_792_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0/$exit
              word_access_0_788_symbol <= Xexit_790_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/word_access_0
            Xexit_787_symbol <= word_access_0_788_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access/$exit
            word_access_785_symbol <= Xexit_787_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/word_access
          Xexit_784_symbol <= word_access_785_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request/$exit
          ptr_deref_215_request_782_symbol <= Xexit_784_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_request
        ptr_deref_215_complete_793: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete 
          signal ptr_deref_215_complete_793_start: Boolean;
          signal Xentry_794_symbol: Boolean;
          signal Xexit_795_symbol: Boolean;
          signal word_access_796_symbol : Boolean;
          signal merge_req_804_symbol : Boolean;
          signal merge_ack_805_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_215_complete_793_start <= ptr_deref_215_active_x_x778_symbol; -- control passed to block
          Xentry_794_symbol  <= ptr_deref_215_complete_793_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/$entry
          word_access_796: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access 
            signal word_access_796_start: Boolean;
            signal Xentry_797_symbol: Boolean;
            signal Xexit_798_symbol: Boolean;
            signal word_access_0_799_symbol : Boolean;
            -- 
          begin -- 
            word_access_796_start <= Xentry_794_symbol; -- control passed to block
            Xentry_797_symbol  <= word_access_796_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/$entry
            word_access_0_799: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0 
              signal word_access_0_799_start: Boolean;
              signal Xentry_800_symbol: Boolean;
              signal Xexit_801_symbol: Boolean;
              signal cr_802_symbol : Boolean;
              signal ca_803_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_799_start <= Xentry_797_symbol; -- control passed to block
              Xentry_800_symbol  <= word_access_0_799_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/$entry
              cr_802_symbol <= Xentry_800_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/cr
              ptr_deref_215_load_0_req_1 <= cr_802_symbol; -- link to DP
              ca_803_symbol <= ptr_deref_215_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/ca
              Xexit_801_symbol <= ca_803_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0/$exit
              word_access_0_799_symbol <= Xexit_801_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/word_access_0
            Xexit_798_symbol <= word_access_0_799_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access/$exit
            word_access_796_symbol <= Xexit_798_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/word_access
          merge_req_804_symbol <= word_access_796_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/merge_req
          ptr_deref_215_gather_scatter_req_0 <= merge_req_804_symbol; -- link to DP
          merge_ack_805_symbol <= ptr_deref_215_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/merge_ack
          Xexit_795_symbol <= merge_ack_805_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete/$exit
          ptr_deref_215_complete_793_symbol <= Xexit_795_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_215_complete
        assign_stmt_221_active_x_x806_symbol <= binary_220_complete_811_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_221_active_
        assign_stmt_221_completed_x_x807_symbol <= assign_stmt_221_active_x_x806_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_221_completed_
        binary_220_active_x_x808_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_active_ 
          signal binary_220_active_x_x808_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_220_active_x_x808_predecessors(0) <= binary_220_trigger_x_x809_symbol;
          binary_220_active_x_x808_predecessors(1) <= simple_obj_ref_218_complete_810_symbol;
          binary_220_active_x_x808_join: join -- 
            port map( -- 
              preds => binary_220_active_x_x808_predecessors,
              symbol_out => binary_220_active_x_x808_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_active_
        binary_220_trigger_x_x809_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_trigger_
        simple_obj_ref_218_complete_810_symbol <= assign_stmt_216_completed_x_x776_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_218_complete
        binary_220_complete_811: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete 
          signal binary_220_complete_811_start: Boolean;
          signal Xentry_812_symbol: Boolean;
          signal Xexit_813_symbol: Boolean;
          signal rr_814_symbol : Boolean;
          signal ra_815_symbol : Boolean;
          signal cr_816_symbol : Boolean;
          signal ca_817_symbol : Boolean;
          -- 
        begin -- 
          binary_220_complete_811_start <= binary_220_active_x_x808_symbol; -- control passed to block
          Xentry_812_symbol  <= binary_220_complete_811_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/$entry
          rr_814_symbol <= Xentry_812_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/rr
          binary_220_inst_req_0 <= rr_814_symbol; -- link to DP
          ra_815_symbol <= binary_220_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/ra
          cr_816_symbol <= ra_815_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/cr
          binary_220_inst_req_1 <= cr_816_symbol; -- link to DP
          ca_817_symbol <= binary_220_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/ca
          Xexit_813_symbol <= ca_817_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete/$exit
          binary_220_complete_811_symbol <= Xexit_813_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/binary_220_complete
        assign_stmt_225_active_x_x818_symbol <= simple_obj_ref_224_complete_820_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_225_active_
        assign_stmt_225_completed_x_x819_symbol <= ptr_deref_223_complete_839_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/assign_stmt_225_completed_
        simple_obj_ref_224_complete_820_symbol <= assign_stmt_221_completed_x_x807_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/simple_obj_ref_224_complete
        ptr_deref_223_trigger_x_x821_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_trigger_ 
          signal ptr_deref_223_trigger_x_x821_predecessors: BooleanArray(4 downto 0);
          -- 
        begin -- 
          ptr_deref_223_trigger_x_x821_predecessors(0) <= ptr_deref_223_word_address_calculated_825_symbol;
          ptr_deref_223_trigger_x_x821_predecessors(1) <= assign_stmt_225_active_x_x818_symbol;
          ptr_deref_223_trigger_x_x821_predecessors(2) <= ptr_deref_183_active_x_x559_symbol;
          ptr_deref_223_trigger_x_x821_predecessors(3) <= ptr_deref_197_active_x_x639_symbol;
          ptr_deref_223_trigger_x_x821_predecessors(4) <= ptr_deref_215_active_x_x778_symbol;
          ptr_deref_223_trigger_x_x821_join: join -- 
            port map( -- 
              preds => ptr_deref_223_trigger_x_x821_predecessors,
              symbol_out => ptr_deref_223_trigger_x_x821_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_trigger_
        ptr_deref_223_active_x_x822_symbol <= ptr_deref_223_request_826_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_active_
        ptr_deref_223_base_address_calculated_823_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_base_address_calculated
        ptr_deref_223_root_address_calculated_824_symbol <= Xentry_554_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_root_address_calculated
        ptr_deref_223_word_address_calculated_825_symbol <= ptr_deref_223_root_address_calculated_824_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_word_address_calculated
        ptr_deref_223_request_826: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request 
          signal ptr_deref_223_request_826_start: Boolean;
          signal Xentry_827_symbol: Boolean;
          signal Xexit_828_symbol: Boolean;
          signal split_req_829_symbol : Boolean;
          signal split_ack_830_symbol : Boolean;
          signal word_access_831_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_223_request_826_start <= ptr_deref_223_trigger_x_x821_symbol; -- control passed to block
          Xentry_827_symbol  <= ptr_deref_223_request_826_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/$entry
          split_req_829_symbol <= Xentry_827_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/split_req
          ptr_deref_223_gather_scatter_req_0 <= split_req_829_symbol; -- link to DP
          split_ack_830_symbol <= ptr_deref_223_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/split_ack
          word_access_831: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access 
            signal word_access_831_start: Boolean;
            signal Xentry_832_symbol: Boolean;
            signal Xexit_833_symbol: Boolean;
            signal word_access_0_834_symbol : Boolean;
            -- 
          begin -- 
            word_access_831_start <= split_ack_830_symbol; -- control passed to block
            Xentry_832_symbol  <= word_access_831_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/$entry
            word_access_0_834: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0 
              signal word_access_0_834_start: Boolean;
              signal Xentry_835_symbol: Boolean;
              signal Xexit_836_symbol: Boolean;
              signal rr_837_symbol : Boolean;
              signal ra_838_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_834_start <= Xentry_832_symbol; -- control passed to block
              Xentry_835_symbol  <= word_access_0_834_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/$entry
              rr_837_symbol <= Xentry_835_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/rr
              ptr_deref_223_store_0_req_0 <= rr_837_symbol; -- link to DP
              ra_838_symbol <= ptr_deref_223_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/ra
              Xexit_836_symbol <= ra_838_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0/$exit
              word_access_0_834_symbol <= Xexit_836_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/word_access_0
            Xexit_833_symbol <= word_access_0_834_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access/$exit
            word_access_831_symbol <= Xexit_833_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/word_access
          Xexit_828_symbol <= word_access_831_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request/$exit
          ptr_deref_223_request_826_symbol <= Xexit_828_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_request
        ptr_deref_223_complete_839: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete 
          signal ptr_deref_223_complete_839_start: Boolean;
          signal Xentry_840_symbol: Boolean;
          signal Xexit_841_symbol: Boolean;
          signal word_access_842_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_223_complete_839_start <= ptr_deref_223_active_x_x822_symbol; -- control passed to block
          Xentry_840_symbol  <= ptr_deref_223_complete_839_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/$entry
          word_access_842: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access 
            signal word_access_842_start: Boolean;
            signal Xentry_843_symbol: Boolean;
            signal Xexit_844_symbol: Boolean;
            signal word_access_0_845_symbol : Boolean;
            -- 
          begin -- 
            word_access_842_start <= Xentry_840_symbol; -- control passed to block
            Xentry_843_symbol  <= word_access_842_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/$entry
            word_access_0_845: Block -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0 
              signal word_access_0_845_start: Boolean;
              signal Xentry_846_symbol: Boolean;
              signal Xexit_847_symbol: Boolean;
              signal cr_848_symbol : Boolean;
              signal ca_849_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_845_start <= Xentry_843_symbol; -- control passed to block
              Xentry_846_symbol  <= word_access_0_845_start; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/$entry
              cr_848_symbol <= Xentry_846_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/cr
              ptr_deref_223_store_0_req_1 <= cr_848_symbol; -- link to DP
              ca_849_symbol <= ptr_deref_223_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/ca
              Xexit_847_symbol <= ca_849_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0/$exit
              word_access_0_845_symbol <= Xexit_847_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/word_access_0
            Xexit_844_symbol <= word_access_0_845_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access/$exit
            word_access_842_symbol <= Xexit_844_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/word_access
          Xexit_841_symbol <= word_access_842_symbol; -- transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete/$exit
          ptr_deref_223_complete_839_symbol <= Xexit_841_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/ptr_deref_223_complete
        Xexit_555_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/$exit 
          signal Xexit_555_predecessors: BooleanArray(5 downto 0);
          -- 
        begin -- 
          Xexit_555_predecessors(0) <= ptr_deref_183_base_address_calculated_560_symbol;
          Xexit_555_predecessors(1) <= ptr_deref_197_base_address_calculated_640_symbol;
          Xexit_555_predecessors(2) <= assign_stmt_212_completed_x_x727_symbol;
          Xexit_555_predecessors(3) <= ptr_deref_215_base_address_calculated_779_symbol;
          Xexit_555_predecessors(4) <= assign_stmt_225_completed_x_x819_symbol;
          Xexit_555_predecessors(5) <= ptr_deref_223_base_address_calculated_823_symbol;
          Xexit_555_join: join -- 
            port map( -- 
              preds => Xexit_555_predecessors,
              symbol_out => Xexit_555_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225/$exit
        assign_stmt_184_to_assign_stmt_225_553_symbol <= Xexit_555_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_184_to_assign_stmt_225
      assign_stmt_233_to_assign_stmt_245_850: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245 
        signal assign_stmt_233_to_assign_stmt_245_850_start: Boolean;
        signal Xentry_851_symbol: Boolean;
        signal Xexit_852_symbol: Boolean;
        signal assign_stmt_237_active_x_x853_symbol : Boolean;
        signal assign_stmt_237_completed_x_x854_symbol : Boolean;
        signal ptr_deref_235_trigger_x_x855_symbol : Boolean;
        signal ptr_deref_235_active_x_x856_symbol : Boolean;
        signal ptr_deref_235_base_address_calculated_857_symbol : Boolean;
        signal ptr_deref_235_root_address_calculated_858_symbol : Boolean;
        signal ptr_deref_235_word_address_calculated_859_symbol : Boolean;
        signal ptr_deref_235_request_860_symbol : Boolean;
        signal ptr_deref_235_complete_873_symbol : Boolean;
        signal assign_stmt_245_active_x_x884_symbol : Boolean;
        signal assign_stmt_245_completed_x_x885_symbol : Boolean;
        signal simple_obj_ref_243_trigger_x_x886_symbol : Boolean;
        signal simple_obj_ref_243_active_x_x887_symbol : Boolean;
        signal simple_obj_ref_243_root_address_calculated_888_symbol : Boolean;
        signal simple_obj_ref_243_word_address_calculated_889_symbol : Boolean;
        signal simple_obj_ref_243_request_890_symbol : Boolean;
        signal simple_obj_ref_243_complete_903_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_233_to_assign_stmt_245_850_start <= assign_stmt_233_to_assign_stmt_245_x_xentry_x_xx_x404_symbol; -- control passed to block
        Xentry_851_symbol  <= assign_stmt_233_to_assign_stmt_245_850_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/$entry
        assign_stmt_237_active_x_x853_symbol <= Xentry_851_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_237_active_
        assign_stmt_237_completed_x_x854_symbol <= ptr_deref_235_complete_873_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_237_completed_
        ptr_deref_235_trigger_x_x855_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_trigger_ 
          signal ptr_deref_235_trigger_x_x855_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_235_trigger_x_x855_predecessors(0) <= ptr_deref_235_word_address_calculated_859_symbol;
          ptr_deref_235_trigger_x_x855_predecessors(1) <= assign_stmt_237_active_x_x853_symbol;
          ptr_deref_235_trigger_x_x855_join: join -- 
            port map( -- 
              preds => ptr_deref_235_trigger_x_x855_predecessors,
              symbol_out => ptr_deref_235_trigger_x_x855_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_trigger_
        ptr_deref_235_active_x_x856_symbol <= ptr_deref_235_request_860_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_active_
        ptr_deref_235_base_address_calculated_857_symbol <= Xentry_851_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_base_address_calculated
        ptr_deref_235_root_address_calculated_858_symbol <= Xentry_851_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_root_address_calculated
        ptr_deref_235_word_address_calculated_859_symbol <= ptr_deref_235_root_address_calculated_858_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_word_address_calculated
        ptr_deref_235_request_860: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request 
          signal ptr_deref_235_request_860_start: Boolean;
          signal Xentry_861_symbol: Boolean;
          signal Xexit_862_symbol: Boolean;
          signal split_req_863_symbol : Boolean;
          signal split_ack_864_symbol : Boolean;
          signal word_access_865_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_235_request_860_start <= ptr_deref_235_trigger_x_x855_symbol; -- control passed to block
          Xentry_861_symbol  <= ptr_deref_235_request_860_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/$entry
          split_req_863_symbol <= Xentry_861_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/split_req
          ptr_deref_235_gather_scatter_req_0 <= split_req_863_symbol; -- link to DP
          split_ack_864_symbol <= ptr_deref_235_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/split_ack
          word_access_865: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access 
            signal word_access_865_start: Boolean;
            signal Xentry_866_symbol: Boolean;
            signal Xexit_867_symbol: Boolean;
            signal word_access_0_868_symbol : Boolean;
            -- 
          begin -- 
            word_access_865_start <= split_ack_864_symbol; -- control passed to block
            Xentry_866_symbol  <= word_access_865_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/$entry
            word_access_0_868: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0 
              signal word_access_0_868_start: Boolean;
              signal Xentry_869_symbol: Boolean;
              signal Xexit_870_symbol: Boolean;
              signal rr_871_symbol : Boolean;
              signal ra_872_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_868_start <= Xentry_866_symbol; -- control passed to block
              Xentry_869_symbol  <= word_access_0_868_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/$entry
              rr_871_symbol <= Xentry_869_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/rr
              ptr_deref_235_store_0_req_0 <= rr_871_symbol; -- link to DP
              ra_872_symbol <= ptr_deref_235_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/ra
              Xexit_870_symbol <= ra_872_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0/$exit
              word_access_0_868_symbol <= Xexit_870_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/word_access_0
            Xexit_867_symbol <= word_access_0_868_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access/$exit
            word_access_865_symbol <= Xexit_867_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/word_access
          Xexit_862_symbol <= word_access_865_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request/$exit
          ptr_deref_235_request_860_symbol <= Xexit_862_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_request
        ptr_deref_235_complete_873: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete 
          signal ptr_deref_235_complete_873_start: Boolean;
          signal Xentry_874_symbol: Boolean;
          signal Xexit_875_symbol: Boolean;
          signal word_access_876_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_235_complete_873_start <= ptr_deref_235_active_x_x856_symbol; -- control passed to block
          Xentry_874_symbol  <= ptr_deref_235_complete_873_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/$entry
          word_access_876: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access 
            signal word_access_876_start: Boolean;
            signal Xentry_877_symbol: Boolean;
            signal Xexit_878_symbol: Boolean;
            signal word_access_0_879_symbol : Boolean;
            -- 
          begin -- 
            word_access_876_start <= Xentry_874_symbol; -- control passed to block
            Xentry_877_symbol  <= word_access_876_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/$entry
            word_access_0_879: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0 
              signal word_access_0_879_start: Boolean;
              signal Xentry_880_symbol: Boolean;
              signal Xexit_881_symbol: Boolean;
              signal cr_882_symbol : Boolean;
              signal ca_883_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_879_start <= Xentry_877_symbol; -- control passed to block
              Xentry_880_symbol  <= word_access_0_879_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/$entry
              cr_882_symbol <= Xentry_880_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/cr
              ptr_deref_235_store_0_req_1 <= cr_882_symbol; -- link to DP
              ca_883_symbol <= ptr_deref_235_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/ca
              Xexit_881_symbol <= ca_883_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0/$exit
              word_access_0_879_symbol <= Xexit_881_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/word_access_0
            Xexit_878_symbol <= word_access_0_879_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access/$exit
            word_access_876_symbol <= Xexit_878_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/word_access
          Xexit_875_symbol <= word_access_876_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete/$exit
          ptr_deref_235_complete_873_symbol <= Xexit_875_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/ptr_deref_235_complete
        assign_stmt_245_active_x_x884_symbol <= Xentry_851_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_245_active_
        assign_stmt_245_completed_x_x885_symbol <= simple_obj_ref_243_complete_903_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/assign_stmt_245_completed_
        simple_obj_ref_243_trigger_x_x886_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_trigger_ 
          signal simple_obj_ref_243_trigger_x_x886_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          simple_obj_ref_243_trigger_x_x886_predecessors(0) <= simple_obj_ref_243_word_address_calculated_889_symbol;
          simple_obj_ref_243_trigger_x_x886_predecessors(1) <= assign_stmt_245_active_x_x884_symbol;
          simple_obj_ref_243_trigger_x_x886_join: join -- 
            port map( -- 
              preds => simple_obj_ref_243_trigger_x_x886_predecessors,
              symbol_out => simple_obj_ref_243_trigger_x_x886_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_trigger_
        simple_obj_ref_243_active_x_x887_symbol <= simple_obj_ref_243_request_890_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_active_
        simple_obj_ref_243_root_address_calculated_888_symbol <= Xentry_851_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_root_address_calculated
        simple_obj_ref_243_word_address_calculated_889_symbol <= simple_obj_ref_243_root_address_calculated_888_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_word_address_calculated
        simple_obj_ref_243_request_890: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request 
          signal simple_obj_ref_243_request_890_start: Boolean;
          signal Xentry_891_symbol: Boolean;
          signal Xexit_892_symbol: Boolean;
          signal split_req_893_symbol : Boolean;
          signal split_ack_894_symbol : Boolean;
          signal word_access_895_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_243_request_890_start <= simple_obj_ref_243_trigger_x_x886_symbol; -- control passed to block
          Xentry_891_symbol  <= simple_obj_ref_243_request_890_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/$entry
          split_req_893_symbol <= Xentry_891_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/split_req
          simple_obj_ref_243_gather_scatter_req_0 <= split_req_893_symbol; -- link to DP
          split_ack_894_symbol <= simple_obj_ref_243_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/split_ack
          word_access_895: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access 
            signal word_access_895_start: Boolean;
            signal Xentry_896_symbol: Boolean;
            signal Xexit_897_symbol: Boolean;
            signal word_access_0_898_symbol : Boolean;
            -- 
          begin -- 
            word_access_895_start <= split_ack_894_symbol; -- control passed to block
            Xentry_896_symbol  <= word_access_895_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/$entry
            word_access_0_898: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0 
              signal word_access_0_898_start: Boolean;
              signal Xentry_899_symbol: Boolean;
              signal Xexit_900_symbol: Boolean;
              signal rr_901_symbol : Boolean;
              signal ra_902_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_898_start <= Xentry_896_symbol; -- control passed to block
              Xentry_899_symbol  <= word_access_0_898_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/$entry
              rr_901_symbol <= Xentry_899_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/rr
              simple_obj_ref_243_store_0_req_0 <= rr_901_symbol; -- link to DP
              ra_902_symbol <= simple_obj_ref_243_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/ra
              Xexit_900_symbol <= ra_902_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0/$exit
              word_access_0_898_symbol <= Xexit_900_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/word_access_0
            Xexit_897_symbol <= word_access_0_898_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access/$exit
            word_access_895_symbol <= Xexit_897_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/word_access
          Xexit_892_symbol <= word_access_895_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request/$exit
          simple_obj_ref_243_request_890_symbol <= Xexit_892_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_request
        simple_obj_ref_243_complete_903: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete 
          signal simple_obj_ref_243_complete_903_start: Boolean;
          signal Xentry_904_symbol: Boolean;
          signal Xexit_905_symbol: Boolean;
          signal word_access_906_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_243_complete_903_start <= simple_obj_ref_243_active_x_x887_symbol; -- control passed to block
          Xentry_904_symbol  <= simple_obj_ref_243_complete_903_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/$entry
          word_access_906: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access 
            signal word_access_906_start: Boolean;
            signal Xentry_907_symbol: Boolean;
            signal Xexit_908_symbol: Boolean;
            signal word_access_0_909_symbol : Boolean;
            -- 
          begin -- 
            word_access_906_start <= Xentry_904_symbol; -- control passed to block
            Xentry_907_symbol  <= word_access_906_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/$entry
            word_access_0_909: Block -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0 
              signal word_access_0_909_start: Boolean;
              signal Xentry_910_symbol: Boolean;
              signal Xexit_911_symbol: Boolean;
              signal cr_912_symbol : Boolean;
              signal ca_913_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_909_start <= Xentry_907_symbol; -- control passed to block
              Xentry_910_symbol  <= word_access_0_909_start; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/$entry
              cr_912_symbol <= Xentry_910_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/cr
              simple_obj_ref_243_store_0_req_1 <= cr_912_symbol; -- link to DP
              ca_913_symbol <= simple_obj_ref_243_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/ca
              Xexit_911_symbol <= ca_913_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0/$exit
              word_access_0_909_symbol <= Xexit_911_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/word_access_0
            Xexit_908_symbol <= word_access_0_909_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access/$exit
            word_access_906_symbol <= Xexit_908_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/word_access
          Xexit_905_symbol <= word_access_906_symbol; -- transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete/$exit
          simple_obj_ref_243_complete_903_symbol <= Xexit_905_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/simple_obj_ref_243_complete
        Xexit_852_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/$exit 
          signal Xexit_852_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          Xexit_852_predecessors(0) <= assign_stmt_237_completed_x_x854_symbol;
          Xexit_852_predecessors(1) <= ptr_deref_235_base_address_calculated_857_symbol;
          Xexit_852_predecessors(2) <= assign_stmt_245_completed_x_x885_symbol;
          Xexit_852_join: join -- 
            port map( -- 
              preds => Xexit_852_predecessors,
              symbol_out => Xexit_852_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245/$exit
        assign_stmt_233_to_assign_stmt_245_850_symbol <= Xexit_852_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_233_to_assign_stmt_245
      assign_stmt_252_914: Block -- branch_block_stmt_134/assign_stmt_252 
        signal assign_stmt_252_914_start: Boolean;
        signal Xentry_915_symbol: Boolean;
        signal Xexit_916_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_252_914_start <= assign_stmt_252_x_xentry_x_xx_x408_symbol; -- control passed to block
        Xentry_915_symbol  <= assign_stmt_252_914_start; -- transition branch_block_stmt_134/assign_stmt_252/$entry
        Xexit_916_symbol <= Xentry_915_symbol; -- transition branch_block_stmt_134/assign_stmt_252/$exit
        assign_stmt_252_914_symbol <= Xexit_916_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_252
      assign_stmt_256_917: Block -- branch_block_stmt_134/assign_stmt_256 
        signal assign_stmt_256_917_start: Boolean;
        signal Xentry_918_symbol: Boolean;
        signal Xexit_919_symbol: Boolean;
        signal assign_stmt_256_active_x_x920_symbol : Boolean;
        signal assign_stmt_256_completed_x_x921_symbol : Boolean;
        signal type_cast_255_active_x_x922_symbol : Boolean;
        signal type_cast_255_trigger_x_x923_symbol : Boolean;
        signal simple_obj_ref_254_trigger_x_x924_symbol : Boolean;
        signal simple_obj_ref_254_complete_925_symbol : Boolean;
        signal type_cast_255_complete_930_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_256_917_start <= assign_stmt_256_x_xentry_x_xx_x410_symbol; -- control passed to block
        Xentry_918_symbol  <= assign_stmt_256_917_start; -- transition branch_block_stmt_134/assign_stmt_256/$entry
        assign_stmt_256_active_x_x920_symbol <= type_cast_255_complete_930_symbol; -- transition branch_block_stmt_134/assign_stmt_256/assign_stmt_256_active_
        assign_stmt_256_completed_x_x921_symbol <= assign_stmt_256_active_x_x920_symbol; -- transition branch_block_stmt_134/assign_stmt_256/assign_stmt_256_completed_
        type_cast_255_active_x_x922_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_256/type_cast_255_active_ 
          signal type_cast_255_active_x_x922_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_255_active_x_x922_predecessors(0) <= type_cast_255_trigger_x_x923_symbol;
          type_cast_255_active_x_x922_predecessors(1) <= simple_obj_ref_254_complete_925_symbol;
          type_cast_255_active_x_x922_join: join -- 
            port map( -- 
              preds => type_cast_255_active_x_x922_predecessors,
              symbol_out => type_cast_255_active_x_x922_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_256/type_cast_255_active_
        type_cast_255_trigger_x_x923_symbol <= Xentry_918_symbol; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_trigger_
        simple_obj_ref_254_trigger_x_x924_symbol <= Xentry_918_symbol; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_trigger_
        simple_obj_ref_254_complete_925: Block -- branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete 
          signal simple_obj_ref_254_complete_925_start: Boolean;
          signal Xentry_926_symbol: Boolean;
          signal Xexit_927_symbol: Boolean;
          signal req_928_symbol : Boolean;
          signal ack_929_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_254_complete_925_start <= simple_obj_ref_254_trigger_x_x924_symbol; -- control passed to block
          Xentry_926_symbol  <= simple_obj_ref_254_complete_925_start; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/$entry
          req_928_symbol <= Xentry_926_symbol; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/req
          simple_obj_ref_254_inst_req_0 <= req_928_symbol; -- link to DP
          ack_929_symbol <= simple_obj_ref_254_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/ack
          Xexit_927_symbol <= ack_929_symbol; -- transition branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete/$exit
          simple_obj_ref_254_complete_925_symbol <= Xexit_927_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_256/simple_obj_ref_254_complete
        type_cast_255_complete_930: Block -- branch_block_stmt_134/assign_stmt_256/type_cast_255_complete 
          signal type_cast_255_complete_930_start: Boolean;
          signal Xentry_931_symbol: Boolean;
          signal Xexit_932_symbol: Boolean;
          signal req_933_symbol : Boolean;
          signal ack_934_symbol : Boolean;
          -- 
        begin -- 
          type_cast_255_complete_930_start <= type_cast_255_active_x_x922_symbol; -- control passed to block
          Xentry_931_symbol  <= type_cast_255_complete_930_start; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/$entry
          req_933_symbol <= Xentry_931_symbol; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/req
          type_cast_255_inst_req_0 <= req_933_symbol; -- link to DP
          ack_934_symbol <= type_cast_255_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/ack
          Xexit_932_symbol <= ack_934_symbol; -- transition branch_block_stmt_134/assign_stmt_256/type_cast_255_complete/$exit
          type_cast_255_complete_930_symbol <= Xexit_932_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_256/type_cast_255_complete
        Xexit_919_symbol <= assign_stmt_256_completed_x_x921_symbol; -- transition branch_block_stmt_134/assign_stmt_256/$exit
        assign_stmt_256_917_symbol <= Xexit_919_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_256
      assign_stmt_260_to_assign_stmt_273_935: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273 
        signal assign_stmt_260_to_assign_stmt_273_935_start: Boolean;
        signal Xentry_936_symbol: Boolean;
        signal Xexit_937_symbol: Boolean;
        signal assign_stmt_260_active_x_x938_symbol : Boolean;
        signal assign_stmt_260_completed_x_x939_symbol : Boolean;
        signal simple_obj_ref_259_complete_940_symbol : Boolean;
        signal ptr_deref_258_trigger_x_x941_symbol : Boolean;
        signal ptr_deref_258_active_x_x942_symbol : Boolean;
        signal ptr_deref_258_base_address_calculated_943_symbol : Boolean;
        signal ptr_deref_258_root_address_calculated_944_symbol : Boolean;
        signal ptr_deref_258_word_address_calculated_945_symbol : Boolean;
        signal ptr_deref_258_request_946_symbol : Boolean;
        signal ptr_deref_258_complete_959_symbol : Boolean;
        signal assign_stmt_264_active_x_x970_symbol : Boolean;
        signal assign_stmt_264_completed_x_x971_symbol : Boolean;
        signal ptr_deref_263_trigger_x_x972_symbol : Boolean;
        signal ptr_deref_263_active_x_x973_symbol : Boolean;
        signal ptr_deref_263_base_address_calculated_974_symbol : Boolean;
        signal ptr_deref_263_root_address_calculated_975_symbol : Boolean;
        signal ptr_deref_263_word_address_calculated_976_symbol : Boolean;
        signal ptr_deref_263_request_977_symbol : Boolean;
        signal ptr_deref_263_complete_988_symbol : Boolean;
        signal assign_stmt_268_active_x_x1001_symbol : Boolean;
        signal assign_stmt_268_completed_x_x1002_symbol : Boolean;
        signal type_cast_267_active_x_x1003_symbol : Boolean;
        signal type_cast_267_trigger_x_x1004_symbol : Boolean;
        signal simple_obj_ref_266_complete_1005_symbol : Boolean;
        signal type_cast_267_complete_1006_symbol : Boolean;
        signal assign_stmt_273_active_x_x1011_symbol : Boolean;
        signal assign_stmt_273_completed_x_x1012_symbol : Boolean;
        signal binary_272_active_x_x1013_symbol : Boolean;
        signal binary_272_trigger_x_x1014_symbol : Boolean;
        signal simple_obj_ref_270_complete_1015_symbol : Boolean;
        signal binary_272_complete_1016_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_260_to_assign_stmt_273_935_start <= assign_stmt_260_to_assign_stmt_273_x_xentry_x_xx_x412_symbol; -- control passed to block
        Xentry_936_symbol  <= assign_stmt_260_to_assign_stmt_273_935_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/$entry
        assign_stmt_260_active_x_x938_symbol <= simple_obj_ref_259_complete_940_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_260_active_
        assign_stmt_260_completed_x_x939_symbol <= ptr_deref_258_complete_959_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_260_completed_
        simple_obj_ref_259_complete_940_symbol <= Xentry_936_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/simple_obj_ref_259_complete
        ptr_deref_258_trigger_x_x941_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_trigger_ 
          signal ptr_deref_258_trigger_x_x941_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_258_trigger_x_x941_predecessors(0) <= ptr_deref_258_word_address_calculated_945_symbol;
          ptr_deref_258_trigger_x_x941_predecessors(1) <= assign_stmt_260_active_x_x938_symbol;
          ptr_deref_258_trigger_x_x941_join: join -- 
            port map( -- 
              preds => ptr_deref_258_trigger_x_x941_predecessors,
              symbol_out => ptr_deref_258_trigger_x_x941_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_trigger_
        ptr_deref_258_active_x_x942_symbol <= ptr_deref_258_request_946_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_active_
        ptr_deref_258_base_address_calculated_943_symbol <= Xentry_936_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_base_address_calculated
        ptr_deref_258_root_address_calculated_944_symbol <= Xentry_936_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_root_address_calculated
        ptr_deref_258_word_address_calculated_945_symbol <= ptr_deref_258_root_address_calculated_944_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_word_address_calculated
        ptr_deref_258_request_946: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request 
          signal ptr_deref_258_request_946_start: Boolean;
          signal Xentry_947_symbol: Boolean;
          signal Xexit_948_symbol: Boolean;
          signal split_req_949_symbol : Boolean;
          signal split_ack_950_symbol : Boolean;
          signal word_access_951_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_258_request_946_start <= ptr_deref_258_trigger_x_x941_symbol; -- control passed to block
          Xentry_947_symbol  <= ptr_deref_258_request_946_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/$entry
          split_req_949_symbol <= Xentry_947_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/split_req
          ptr_deref_258_gather_scatter_req_0 <= split_req_949_symbol; -- link to DP
          split_ack_950_symbol <= ptr_deref_258_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/split_ack
          word_access_951: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access 
            signal word_access_951_start: Boolean;
            signal Xentry_952_symbol: Boolean;
            signal Xexit_953_symbol: Boolean;
            signal word_access_0_954_symbol : Boolean;
            -- 
          begin -- 
            word_access_951_start <= split_ack_950_symbol; -- control passed to block
            Xentry_952_symbol  <= word_access_951_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/$entry
            word_access_0_954: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0 
              signal word_access_0_954_start: Boolean;
              signal Xentry_955_symbol: Boolean;
              signal Xexit_956_symbol: Boolean;
              signal rr_957_symbol : Boolean;
              signal ra_958_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_954_start <= Xentry_952_symbol; -- control passed to block
              Xentry_955_symbol  <= word_access_0_954_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/$entry
              rr_957_symbol <= Xentry_955_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/rr
              ptr_deref_258_store_0_req_0 <= rr_957_symbol; -- link to DP
              ra_958_symbol <= ptr_deref_258_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/ra
              Xexit_956_symbol <= ra_958_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0/$exit
              word_access_0_954_symbol <= Xexit_956_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/word_access_0
            Xexit_953_symbol <= word_access_0_954_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access/$exit
            word_access_951_symbol <= Xexit_953_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/word_access
          Xexit_948_symbol <= word_access_951_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request/$exit
          ptr_deref_258_request_946_symbol <= Xexit_948_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_request
        ptr_deref_258_complete_959: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete 
          signal ptr_deref_258_complete_959_start: Boolean;
          signal Xentry_960_symbol: Boolean;
          signal Xexit_961_symbol: Boolean;
          signal word_access_962_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_258_complete_959_start <= ptr_deref_258_active_x_x942_symbol; -- control passed to block
          Xentry_960_symbol  <= ptr_deref_258_complete_959_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/$entry
          word_access_962: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access 
            signal word_access_962_start: Boolean;
            signal Xentry_963_symbol: Boolean;
            signal Xexit_964_symbol: Boolean;
            signal word_access_0_965_symbol : Boolean;
            -- 
          begin -- 
            word_access_962_start <= Xentry_960_symbol; -- control passed to block
            Xentry_963_symbol  <= word_access_962_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/$entry
            word_access_0_965: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0 
              signal word_access_0_965_start: Boolean;
              signal Xentry_966_symbol: Boolean;
              signal Xexit_967_symbol: Boolean;
              signal cr_968_symbol : Boolean;
              signal ca_969_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_965_start <= Xentry_963_symbol; -- control passed to block
              Xentry_966_symbol  <= word_access_0_965_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/$entry
              cr_968_symbol <= Xentry_966_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/cr
              ptr_deref_258_store_0_req_1 <= cr_968_symbol; -- link to DP
              ca_969_symbol <= ptr_deref_258_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/ca
              Xexit_967_symbol <= ca_969_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0/$exit
              word_access_0_965_symbol <= Xexit_967_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/word_access_0
            Xexit_964_symbol <= word_access_0_965_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access/$exit
            word_access_962_symbol <= Xexit_964_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/word_access
          Xexit_961_symbol <= word_access_962_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete/$exit
          ptr_deref_258_complete_959_symbol <= Xexit_961_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_258_complete
        assign_stmt_264_active_x_x970_symbol <= ptr_deref_263_complete_988_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_264_active_
        assign_stmt_264_completed_x_x971_symbol <= assign_stmt_264_active_x_x970_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_264_completed_
        ptr_deref_263_trigger_x_x972_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_trigger_ 
          signal ptr_deref_263_trigger_x_x972_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_263_trigger_x_x972_predecessors(0) <= ptr_deref_263_word_address_calculated_976_symbol;
          ptr_deref_263_trigger_x_x972_predecessors(1) <= ptr_deref_258_active_x_x942_symbol;
          ptr_deref_263_trigger_x_x972_join: join -- 
            port map( -- 
              preds => ptr_deref_263_trigger_x_x972_predecessors,
              symbol_out => ptr_deref_263_trigger_x_x972_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_trigger_
        ptr_deref_263_active_x_x973_symbol <= ptr_deref_263_request_977_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_active_
        ptr_deref_263_base_address_calculated_974_symbol <= Xentry_936_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_base_address_calculated
        ptr_deref_263_root_address_calculated_975_symbol <= Xentry_936_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_root_address_calculated
        ptr_deref_263_word_address_calculated_976_symbol <= ptr_deref_263_root_address_calculated_975_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_word_address_calculated
        ptr_deref_263_request_977: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request 
          signal ptr_deref_263_request_977_start: Boolean;
          signal Xentry_978_symbol: Boolean;
          signal Xexit_979_symbol: Boolean;
          signal word_access_980_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_263_request_977_start <= ptr_deref_263_trigger_x_x972_symbol; -- control passed to block
          Xentry_978_symbol  <= ptr_deref_263_request_977_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/$entry
          word_access_980: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access 
            signal word_access_980_start: Boolean;
            signal Xentry_981_symbol: Boolean;
            signal Xexit_982_symbol: Boolean;
            signal word_access_0_983_symbol : Boolean;
            -- 
          begin -- 
            word_access_980_start <= Xentry_978_symbol; -- control passed to block
            Xentry_981_symbol  <= word_access_980_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/$entry
            word_access_0_983: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0 
              signal word_access_0_983_start: Boolean;
              signal Xentry_984_symbol: Boolean;
              signal Xexit_985_symbol: Boolean;
              signal rr_986_symbol : Boolean;
              signal ra_987_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_983_start <= Xentry_981_symbol; -- control passed to block
              Xentry_984_symbol  <= word_access_0_983_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/$entry
              rr_986_symbol <= Xentry_984_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/rr
              ptr_deref_263_load_0_req_0 <= rr_986_symbol; -- link to DP
              ra_987_symbol <= ptr_deref_263_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/ra
              Xexit_985_symbol <= ra_987_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0/$exit
              word_access_0_983_symbol <= Xexit_985_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/word_access_0
            Xexit_982_symbol <= word_access_0_983_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access/$exit
            word_access_980_symbol <= Xexit_982_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/word_access
          Xexit_979_symbol <= word_access_980_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request/$exit
          ptr_deref_263_request_977_symbol <= Xexit_979_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_request
        ptr_deref_263_complete_988: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete 
          signal ptr_deref_263_complete_988_start: Boolean;
          signal Xentry_989_symbol: Boolean;
          signal Xexit_990_symbol: Boolean;
          signal word_access_991_symbol : Boolean;
          signal merge_req_999_symbol : Boolean;
          signal merge_ack_1000_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_263_complete_988_start <= ptr_deref_263_active_x_x973_symbol; -- control passed to block
          Xentry_989_symbol  <= ptr_deref_263_complete_988_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/$entry
          word_access_991: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access 
            signal word_access_991_start: Boolean;
            signal Xentry_992_symbol: Boolean;
            signal Xexit_993_symbol: Boolean;
            signal word_access_0_994_symbol : Boolean;
            -- 
          begin -- 
            word_access_991_start <= Xentry_989_symbol; -- control passed to block
            Xentry_992_symbol  <= word_access_991_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/$entry
            word_access_0_994: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0 
              signal word_access_0_994_start: Boolean;
              signal Xentry_995_symbol: Boolean;
              signal Xexit_996_symbol: Boolean;
              signal cr_997_symbol : Boolean;
              signal ca_998_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_994_start <= Xentry_992_symbol; -- control passed to block
              Xentry_995_symbol  <= word_access_0_994_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/$entry
              cr_997_symbol <= Xentry_995_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/cr
              ptr_deref_263_load_0_req_1 <= cr_997_symbol; -- link to DP
              ca_998_symbol <= ptr_deref_263_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/ca
              Xexit_996_symbol <= ca_998_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0/$exit
              word_access_0_994_symbol <= Xexit_996_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/word_access_0
            Xexit_993_symbol <= word_access_0_994_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access/$exit
            word_access_991_symbol <= Xexit_993_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/word_access
          merge_req_999_symbol <= word_access_991_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/merge_req
          ptr_deref_263_gather_scatter_req_0 <= merge_req_999_symbol; -- link to DP
          merge_ack_1000_symbol <= ptr_deref_263_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/merge_ack
          Xexit_990_symbol <= merge_ack_1000_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete/$exit
          ptr_deref_263_complete_988_symbol <= Xexit_990_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/ptr_deref_263_complete
        assign_stmt_268_active_x_x1001_symbol <= type_cast_267_complete_1006_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_268_active_
        assign_stmt_268_completed_x_x1002_symbol <= assign_stmt_268_active_x_x1001_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_268_completed_
        type_cast_267_active_x_x1003_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_active_ 
          signal type_cast_267_active_x_x1003_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_267_active_x_x1003_predecessors(0) <= type_cast_267_trigger_x_x1004_symbol;
          type_cast_267_active_x_x1003_predecessors(1) <= simple_obj_ref_266_complete_1005_symbol;
          type_cast_267_active_x_x1003_join: join -- 
            port map( -- 
              preds => type_cast_267_active_x_x1003_predecessors,
              symbol_out => type_cast_267_active_x_x1003_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_active_
        type_cast_267_trigger_x_x1004_symbol <= Xentry_936_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_trigger_
        simple_obj_ref_266_complete_1005_symbol <= assign_stmt_264_completed_x_x971_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/simple_obj_ref_266_complete
        type_cast_267_complete_1006: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete 
          signal type_cast_267_complete_1006_start: Boolean;
          signal Xentry_1007_symbol: Boolean;
          signal Xexit_1008_symbol: Boolean;
          signal req_1009_symbol : Boolean;
          signal ack_1010_symbol : Boolean;
          -- 
        begin -- 
          type_cast_267_complete_1006_start <= type_cast_267_active_x_x1003_symbol; -- control passed to block
          Xentry_1007_symbol  <= type_cast_267_complete_1006_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/$entry
          req_1009_symbol <= Xentry_1007_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/req
          type_cast_267_inst_req_0 <= req_1009_symbol; -- link to DP
          ack_1010_symbol <= type_cast_267_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/ack
          Xexit_1008_symbol <= ack_1010_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete/$exit
          type_cast_267_complete_1006_symbol <= Xexit_1008_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/type_cast_267_complete
        assign_stmt_273_active_x_x1011_symbol <= binary_272_complete_1016_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_273_active_
        assign_stmt_273_completed_x_x1012_symbol <= assign_stmt_273_active_x_x1011_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/assign_stmt_273_completed_
        binary_272_active_x_x1013_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_active_ 
          signal binary_272_active_x_x1013_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_272_active_x_x1013_predecessors(0) <= binary_272_trigger_x_x1014_symbol;
          binary_272_active_x_x1013_predecessors(1) <= simple_obj_ref_270_complete_1015_symbol;
          binary_272_active_x_x1013_join: join -- 
            port map( -- 
              preds => binary_272_active_x_x1013_predecessors,
              symbol_out => binary_272_active_x_x1013_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_active_
        binary_272_trigger_x_x1014_symbol <= Xentry_936_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_trigger_
        simple_obj_ref_270_complete_1015_symbol <= assign_stmt_268_completed_x_x1002_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/simple_obj_ref_270_complete
        binary_272_complete_1016: Block -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete 
          signal binary_272_complete_1016_start: Boolean;
          signal Xentry_1017_symbol: Boolean;
          signal Xexit_1018_symbol: Boolean;
          signal rr_1019_symbol : Boolean;
          signal ra_1020_symbol : Boolean;
          signal cr_1021_symbol : Boolean;
          signal ca_1022_symbol : Boolean;
          -- 
        begin -- 
          binary_272_complete_1016_start <= binary_272_active_x_x1013_symbol; -- control passed to block
          Xentry_1017_symbol  <= binary_272_complete_1016_start; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/$entry
          rr_1019_symbol <= Xentry_1017_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/rr
          binary_272_inst_req_0 <= rr_1019_symbol; -- link to DP
          ra_1020_symbol <= binary_272_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/ra
          cr_1021_symbol <= ra_1020_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/cr
          binary_272_inst_req_1 <= cr_1021_symbol; -- link to DP
          ca_1022_symbol <= binary_272_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/ca
          Xexit_1018_symbol <= ca_1022_symbol; -- transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete/$exit
          binary_272_complete_1016_symbol <= Xexit_1018_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/binary_272_complete
        Xexit_937_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/$exit 
          signal Xexit_937_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          Xexit_937_predecessors(0) <= assign_stmt_260_completed_x_x939_symbol;
          Xexit_937_predecessors(1) <= ptr_deref_258_base_address_calculated_943_symbol;
          Xexit_937_predecessors(2) <= ptr_deref_263_base_address_calculated_974_symbol;
          Xexit_937_predecessors(3) <= assign_stmt_273_completed_x_x1012_symbol;
          Xexit_937_join: join -- 
            port map( -- 
              preds => Xexit_937_predecessors,
              symbol_out => Xexit_937_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273/$exit
        assign_stmt_260_to_assign_stmt_273_935_symbol <= Xexit_937_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_260_to_assign_stmt_273
      if_stmt_274_dead_link_1023: Block -- branch_block_stmt_134/if_stmt_274_dead_link 
        signal if_stmt_274_dead_link_1023_start: Boolean;
        signal Xentry_1024_symbol: Boolean;
        signal Xexit_1025_symbol: Boolean;
        signal dead_transition_1026_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_dead_link_1023_start <= if_stmt_274_x_xentry_x_xx_x414_symbol; -- control passed to block
        Xentry_1024_symbol  <= if_stmt_274_dead_link_1023_start; -- transition branch_block_stmt_134/if_stmt_274_dead_link/$entry
        dead_transition_1026_symbol <= false;
        Xexit_1025_symbol <= dead_transition_1026_symbol; -- transition branch_block_stmt_134/if_stmt_274_dead_link/$exit
        if_stmt_274_dead_link_1023_symbol <= Xexit_1025_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_dead_link
      if_stmt_274_eval_test_1027: Block -- branch_block_stmt_134/if_stmt_274_eval_test 
        signal if_stmt_274_eval_test_1027_start: Boolean;
        signal Xentry_1028_symbol: Boolean;
        signal Xexit_1029_symbol: Boolean;
        signal branch_req_1030_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_eval_test_1027_start <= if_stmt_274_x_xentry_x_xx_x414_symbol; -- control passed to block
        Xentry_1028_symbol  <= if_stmt_274_eval_test_1027_start; -- transition branch_block_stmt_134/if_stmt_274_eval_test/$entry
        branch_req_1030_symbol <= Xentry_1028_symbol; -- transition branch_block_stmt_134/if_stmt_274_eval_test/branch_req
        if_stmt_274_branch_req_0 <= branch_req_1030_symbol; -- link to DP
        Xexit_1029_symbol <= branch_req_1030_symbol; -- transition branch_block_stmt_134/if_stmt_274_eval_test/$exit
        if_stmt_274_eval_test_1027_symbol <= Xexit_1029_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_eval_test
      simple_obj_ref_275_place_1031_symbol  <=  if_stmt_274_eval_test_1027_symbol; -- place branch_block_stmt_134/simple_obj_ref_275_place (optimized away) 
      if_stmt_274_if_link_1032: Block -- branch_block_stmt_134/if_stmt_274_if_link 
        signal if_stmt_274_if_link_1032_start: Boolean;
        signal Xentry_1033_symbol: Boolean;
        signal Xexit_1034_symbol: Boolean;
        signal if_choice_transition_1035_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_if_link_1032_start <= simple_obj_ref_275_place_1031_symbol; -- control passed to block
        Xentry_1033_symbol  <= if_stmt_274_if_link_1032_start; -- transition branch_block_stmt_134/if_stmt_274_if_link/$entry
        if_choice_transition_1035_symbol <= if_stmt_274_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_274_if_link/if_choice_transition
        Xexit_1034_symbol <= if_choice_transition_1035_symbol; -- transition branch_block_stmt_134/if_stmt_274_if_link/$exit
        if_stmt_274_if_link_1032_symbol <= Xexit_1034_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_if_link
      if_stmt_274_else_link_1036: Block -- branch_block_stmt_134/if_stmt_274_else_link 
        signal if_stmt_274_else_link_1036_start: Boolean;
        signal Xentry_1037_symbol: Boolean;
        signal Xexit_1038_symbol: Boolean;
        signal else_choice_transition_1039_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_274_else_link_1036_start <= simple_obj_ref_275_place_1031_symbol; -- control passed to block
        Xentry_1037_symbol  <= if_stmt_274_else_link_1036_start; -- transition branch_block_stmt_134/if_stmt_274_else_link/$entry
        else_choice_transition_1039_symbol <= if_stmt_274_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_274_else_link/else_choice_transition
        Xexit_1038_symbol <= else_choice_transition_1039_symbol; -- transition branch_block_stmt_134/if_stmt_274_else_link/$exit
        if_stmt_274_else_link_1036_symbol <= Xexit_1038_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_274_else_link
      bb_4_bb_5_1040_symbol  <=  if_stmt_274_if_link_1032_symbol; -- place branch_block_stmt_134/bb_4_bb_5 (optimized away) 
      bb_4_bb_8_1041_symbol  <=  if_stmt_274_else_link_1036_symbol; -- place branch_block_stmt_134/bb_4_bb_8 (optimized away) 
      assign_stmt_283_to_assign_stmt_297_1042: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297 
        signal assign_stmt_283_to_assign_stmt_297_1042_start: Boolean;
        signal Xentry_1043_symbol: Boolean;
        signal Xexit_1044_symbol: Boolean;
        signal assign_stmt_283_active_x_x1045_symbol : Boolean;
        signal assign_stmt_283_completed_x_x1046_symbol : Boolean;
        signal simple_obj_ref_282_trigger_x_x1047_symbol : Boolean;
        signal simple_obj_ref_282_active_x_x1048_symbol : Boolean;
        signal simple_obj_ref_282_root_address_calculated_1049_symbol : Boolean;
        signal simple_obj_ref_282_word_address_calculated_1050_symbol : Boolean;
        signal simple_obj_ref_282_request_1051_symbol : Boolean;
        signal simple_obj_ref_282_complete_1062_symbol : Boolean;
        signal assign_stmt_287_active_x_x1075_symbol : Boolean;
        signal assign_stmt_287_completed_x_x1076_symbol : Boolean;
        signal simple_obj_ref_286_complete_1077_symbol : Boolean;
        signal ptr_deref_285_trigger_x_x1078_symbol : Boolean;
        signal ptr_deref_285_active_x_x1079_symbol : Boolean;
        signal ptr_deref_285_base_address_calculated_1080_symbol : Boolean;
        signal ptr_deref_285_root_address_calculated_1081_symbol : Boolean;
        signal ptr_deref_285_word_address_calculated_1082_symbol : Boolean;
        signal ptr_deref_285_request_1083_symbol : Boolean;
        signal ptr_deref_285_complete_1096_symbol : Boolean;
        signal assign_stmt_290_active_x_x1107_symbol : Boolean;
        signal assign_stmt_290_completed_x_x1108_symbol : Boolean;
        signal simple_obj_ref_289_trigger_x_x1109_symbol : Boolean;
        signal simple_obj_ref_289_active_x_x1110_symbol : Boolean;
        signal simple_obj_ref_289_root_address_calculated_1111_symbol : Boolean;
        signal simple_obj_ref_289_word_address_calculated_1112_symbol : Boolean;
        signal simple_obj_ref_289_request_1113_symbol : Boolean;
        signal simple_obj_ref_289_complete_1124_symbol : Boolean;
        signal assign_stmt_297_active_x_x1137_symbol : Boolean;
        signal assign_stmt_297_completed_x_x1138_symbol : Boolean;
        signal binary_296_active_x_x1139_symbol : Boolean;
        signal binary_296_trigger_x_x1140_symbol : Boolean;
        signal type_cast_293_active_x_x1141_symbol : Boolean;
        signal type_cast_293_trigger_x_x1142_symbol : Boolean;
        signal simple_obj_ref_292_complete_1143_symbol : Boolean;
        signal type_cast_293_complete_1144_symbol : Boolean;
        signal binary_296_complete_1149_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_283_to_assign_stmt_297_1042_start <= assign_stmt_283_to_assign_stmt_297_x_xentry_x_xx_x418_symbol; -- control passed to block
        Xentry_1043_symbol  <= assign_stmt_283_to_assign_stmt_297_1042_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/$entry
        assign_stmt_283_active_x_x1045_symbol <= simple_obj_ref_282_complete_1062_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_283_active_
        assign_stmt_283_completed_x_x1046_symbol <= assign_stmt_283_active_x_x1045_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_283_completed_
        simple_obj_ref_282_trigger_x_x1047_symbol <= simple_obj_ref_282_word_address_calculated_1050_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_trigger_
        simple_obj_ref_282_active_x_x1048_symbol <= simple_obj_ref_282_request_1051_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_active_
        simple_obj_ref_282_root_address_calculated_1049_symbol <= Xentry_1043_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_root_address_calculated
        simple_obj_ref_282_word_address_calculated_1050_symbol <= simple_obj_ref_282_root_address_calculated_1049_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_word_address_calculated
        simple_obj_ref_282_request_1051: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request 
          signal simple_obj_ref_282_request_1051_start: Boolean;
          signal Xentry_1052_symbol: Boolean;
          signal Xexit_1053_symbol: Boolean;
          signal word_access_1054_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_282_request_1051_start <= simple_obj_ref_282_trigger_x_x1047_symbol; -- control passed to block
          Xentry_1052_symbol  <= simple_obj_ref_282_request_1051_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/$entry
          word_access_1054: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access 
            signal word_access_1054_start: Boolean;
            signal Xentry_1055_symbol: Boolean;
            signal Xexit_1056_symbol: Boolean;
            signal word_access_0_1057_symbol : Boolean;
            -- 
          begin -- 
            word_access_1054_start <= Xentry_1052_symbol; -- control passed to block
            Xentry_1055_symbol  <= word_access_1054_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/$entry
            word_access_0_1057: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0 
              signal word_access_0_1057_start: Boolean;
              signal Xentry_1058_symbol: Boolean;
              signal Xexit_1059_symbol: Boolean;
              signal rr_1060_symbol : Boolean;
              signal ra_1061_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1057_start <= Xentry_1055_symbol; -- control passed to block
              Xentry_1058_symbol  <= word_access_0_1057_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/$entry
              rr_1060_symbol <= Xentry_1058_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/rr
              simple_obj_ref_282_load_0_req_0 <= rr_1060_symbol; -- link to DP
              ra_1061_symbol <= simple_obj_ref_282_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/ra
              Xexit_1059_symbol <= ra_1061_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0/$exit
              word_access_0_1057_symbol <= Xexit_1059_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/word_access_0
            Xexit_1056_symbol <= word_access_0_1057_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access/$exit
            word_access_1054_symbol <= Xexit_1056_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/word_access
          Xexit_1053_symbol <= word_access_1054_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request/$exit
          simple_obj_ref_282_request_1051_symbol <= Xexit_1053_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_request
        simple_obj_ref_282_complete_1062: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete 
          signal simple_obj_ref_282_complete_1062_start: Boolean;
          signal Xentry_1063_symbol: Boolean;
          signal Xexit_1064_symbol: Boolean;
          signal word_access_1065_symbol : Boolean;
          signal merge_req_1073_symbol : Boolean;
          signal merge_ack_1074_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_282_complete_1062_start <= simple_obj_ref_282_active_x_x1048_symbol; -- control passed to block
          Xentry_1063_symbol  <= simple_obj_ref_282_complete_1062_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/$entry
          word_access_1065: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access 
            signal word_access_1065_start: Boolean;
            signal Xentry_1066_symbol: Boolean;
            signal Xexit_1067_symbol: Boolean;
            signal word_access_0_1068_symbol : Boolean;
            -- 
          begin -- 
            word_access_1065_start <= Xentry_1063_symbol; -- control passed to block
            Xentry_1066_symbol  <= word_access_1065_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/$entry
            word_access_0_1068: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0 
              signal word_access_0_1068_start: Boolean;
              signal Xentry_1069_symbol: Boolean;
              signal Xexit_1070_symbol: Boolean;
              signal cr_1071_symbol : Boolean;
              signal ca_1072_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1068_start <= Xentry_1066_symbol; -- control passed to block
              Xentry_1069_symbol  <= word_access_0_1068_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/$entry
              cr_1071_symbol <= Xentry_1069_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/cr
              simple_obj_ref_282_load_0_req_1 <= cr_1071_symbol; -- link to DP
              ca_1072_symbol <= simple_obj_ref_282_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/ca
              Xexit_1070_symbol <= ca_1072_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0/$exit
              word_access_0_1068_symbol <= Xexit_1070_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/word_access_0
            Xexit_1067_symbol <= word_access_0_1068_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access/$exit
            word_access_1065_symbol <= Xexit_1067_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/word_access
          merge_req_1073_symbol <= word_access_1065_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/merge_req
          simple_obj_ref_282_gather_scatter_req_0 <= merge_req_1073_symbol; -- link to DP
          merge_ack_1074_symbol <= simple_obj_ref_282_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/merge_ack
          Xexit_1064_symbol <= merge_ack_1074_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete/$exit
          simple_obj_ref_282_complete_1062_symbol <= Xexit_1064_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_282_complete
        assign_stmt_287_active_x_x1075_symbol <= simple_obj_ref_286_complete_1077_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_287_active_
        assign_stmt_287_completed_x_x1076_symbol <= ptr_deref_285_complete_1096_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_287_completed_
        simple_obj_ref_286_complete_1077_symbol <= assign_stmt_283_completed_x_x1046_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_286_complete
        ptr_deref_285_trigger_x_x1078_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_trigger_ 
          signal ptr_deref_285_trigger_x_x1078_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_285_trigger_x_x1078_predecessors(0) <= ptr_deref_285_word_address_calculated_1082_symbol;
          ptr_deref_285_trigger_x_x1078_predecessors(1) <= assign_stmt_287_active_x_x1075_symbol;
          ptr_deref_285_trigger_x_x1078_join: join -- 
            port map( -- 
              preds => ptr_deref_285_trigger_x_x1078_predecessors,
              symbol_out => ptr_deref_285_trigger_x_x1078_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_trigger_
        ptr_deref_285_active_x_x1079_symbol <= ptr_deref_285_request_1083_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_active_
        ptr_deref_285_base_address_calculated_1080_symbol <= Xentry_1043_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_base_address_calculated
        ptr_deref_285_root_address_calculated_1081_symbol <= Xentry_1043_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_root_address_calculated
        ptr_deref_285_word_address_calculated_1082_symbol <= ptr_deref_285_root_address_calculated_1081_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_word_address_calculated
        ptr_deref_285_request_1083: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request 
          signal ptr_deref_285_request_1083_start: Boolean;
          signal Xentry_1084_symbol: Boolean;
          signal Xexit_1085_symbol: Boolean;
          signal split_req_1086_symbol : Boolean;
          signal split_ack_1087_symbol : Boolean;
          signal word_access_1088_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_285_request_1083_start <= ptr_deref_285_trigger_x_x1078_symbol; -- control passed to block
          Xentry_1084_symbol  <= ptr_deref_285_request_1083_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/$entry
          split_req_1086_symbol <= Xentry_1084_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/split_req
          ptr_deref_285_gather_scatter_req_0 <= split_req_1086_symbol; -- link to DP
          split_ack_1087_symbol <= ptr_deref_285_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/split_ack
          word_access_1088: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access 
            signal word_access_1088_start: Boolean;
            signal Xentry_1089_symbol: Boolean;
            signal Xexit_1090_symbol: Boolean;
            signal word_access_0_1091_symbol : Boolean;
            -- 
          begin -- 
            word_access_1088_start <= split_ack_1087_symbol; -- control passed to block
            Xentry_1089_symbol  <= word_access_1088_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/$entry
            word_access_0_1091: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0 
              signal word_access_0_1091_start: Boolean;
              signal Xentry_1092_symbol: Boolean;
              signal Xexit_1093_symbol: Boolean;
              signal rr_1094_symbol : Boolean;
              signal ra_1095_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1091_start <= Xentry_1089_symbol; -- control passed to block
              Xentry_1092_symbol  <= word_access_0_1091_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/$entry
              rr_1094_symbol <= Xentry_1092_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/rr
              ptr_deref_285_store_0_req_0 <= rr_1094_symbol; -- link to DP
              ra_1095_symbol <= ptr_deref_285_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/ra
              Xexit_1093_symbol <= ra_1095_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0/$exit
              word_access_0_1091_symbol <= Xexit_1093_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/word_access_0
            Xexit_1090_symbol <= word_access_0_1091_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access/$exit
            word_access_1088_symbol <= Xexit_1090_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/word_access
          Xexit_1085_symbol <= word_access_1088_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request/$exit
          ptr_deref_285_request_1083_symbol <= Xexit_1085_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_request
        ptr_deref_285_complete_1096: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete 
          signal ptr_deref_285_complete_1096_start: Boolean;
          signal Xentry_1097_symbol: Boolean;
          signal Xexit_1098_symbol: Boolean;
          signal word_access_1099_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_285_complete_1096_start <= ptr_deref_285_active_x_x1079_symbol; -- control passed to block
          Xentry_1097_symbol  <= ptr_deref_285_complete_1096_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/$entry
          word_access_1099: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access 
            signal word_access_1099_start: Boolean;
            signal Xentry_1100_symbol: Boolean;
            signal Xexit_1101_symbol: Boolean;
            signal word_access_0_1102_symbol : Boolean;
            -- 
          begin -- 
            word_access_1099_start <= Xentry_1097_symbol; -- control passed to block
            Xentry_1100_symbol  <= word_access_1099_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/$entry
            word_access_0_1102: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0 
              signal word_access_0_1102_start: Boolean;
              signal Xentry_1103_symbol: Boolean;
              signal Xexit_1104_symbol: Boolean;
              signal cr_1105_symbol : Boolean;
              signal ca_1106_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1102_start <= Xentry_1100_symbol; -- control passed to block
              Xentry_1103_symbol  <= word_access_0_1102_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/$entry
              cr_1105_symbol <= Xentry_1103_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/cr
              ptr_deref_285_store_0_req_1 <= cr_1105_symbol; -- link to DP
              ca_1106_symbol <= ptr_deref_285_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/ca
              Xexit_1104_symbol <= ca_1106_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0/$exit
              word_access_0_1102_symbol <= Xexit_1104_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/word_access_0
            Xexit_1101_symbol <= word_access_0_1102_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access/$exit
            word_access_1099_symbol <= Xexit_1101_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/word_access
          Xexit_1098_symbol <= word_access_1099_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete/$exit
          ptr_deref_285_complete_1096_symbol <= Xexit_1098_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/ptr_deref_285_complete
        assign_stmt_290_active_x_x1107_symbol <= simple_obj_ref_289_complete_1124_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_290_active_
        assign_stmt_290_completed_x_x1108_symbol <= assign_stmt_290_active_x_x1107_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_290_completed_
        simple_obj_ref_289_trigger_x_x1109_symbol <= simple_obj_ref_289_word_address_calculated_1112_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_trigger_
        simple_obj_ref_289_active_x_x1110_symbol <= simple_obj_ref_289_request_1113_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_active_
        simple_obj_ref_289_root_address_calculated_1111_symbol <= Xentry_1043_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_root_address_calculated
        simple_obj_ref_289_word_address_calculated_1112_symbol <= simple_obj_ref_289_root_address_calculated_1111_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_word_address_calculated
        simple_obj_ref_289_request_1113: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request 
          signal simple_obj_ref_289_request_1113_start: Boolean;
          signal Xentry_1114_symbol: Boolean;
          signal Xexit_1115_symbol: Boolean;
          signal word_access_1116_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_289_request_1113_start <= simple_obj_ref_289_trigger_x_x1109_symbol; -- control passed to block
          Xentry_1114_symbol  <= simple_obj_ref_289_request_1113_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/$entry
          word_access_1116: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access 
            signal word_access_1116_start: Boolean;
            signal Xentry_1117_symbol: Boolean;
            signal Xexit_1118_symbol: Boolean;
            signal word_access_0_1119_symbol : Boolean;
            -- 
          begin -- 
            word_access_1116_start <= Xentry_1114_symbol; -- control passed to block
            Xentry_1117_symbol  <= word_access_1116_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/$entry
            word_access_0_1119: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0 
              signal word_access_0_1119_start: Boolean;
              signal Xentry_1120_symbol: Boolean;
              signal Xexit_1121_symbol: Boolean;
              signal rr_1122_symbol : Boolean;
              signal ra_1123_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1119_start <= Xentry_1117_symbol; -- control passed to block
              Xentry_1120_symbol  <= word_access_0_1119_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/$entry
              rr_1122_symbol <= Xentry_1120_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/rr
              simple_obj_ref_289_load_0_req_0 <= rr_1122_symbol; -- link to DP
              ra_1123_symbol <= simple_obj_ref_289_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/ra
              Xexit_1121_symbol <= ra_1123_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0/$exit
              word_access_0_1119_symbol <= Xexit_1121_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/word_access_0
            Xexit_1118_symbol <= word_access_0_1119_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access/$exit
            word_access_1116_symbol <= Xexit_1118_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/word_access
          Xexit_1115_symbol <= word_access_1116_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request/$exit
          simple_obj_ref_289_request_1113_symbol <= Xexit_1115_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_request
        simple_obj_ref_289_complete_1124: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete 
          signal simple_obj_ref_289_complete_1124_start: Boolean;
          signal Xentry_1125_symbol: Boolean;
          signal Xexit_1126_symbol: Boolean;
          signal word_access_1127_symbol : Boolean;
          signal merge_req_1135_symbol : Boolean;
          signal merge_ack_1136_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_289_complete_1124_start <= simple_obj_ref_289_active_x_x1110_symbol; -- control passed to block
          Xentry_1125_symbol  <= simple_obj_ref_289_complete_1124_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/$entry
          word_access_1127: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access 
            signal word_access_1127_start: Boolean;
            signal Xentry_1128_symbol: Boolean;
            signal Xexit_1129_symbol: Boolean;
            signal word_access_0_1130_symbol : Boolean;
            -- 
          begin -- 
            word_access_1127_start <= Xentry_1125_symbol; -- control passed to block
            Xentry_1128_symbol  <= word_access_1127_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/$entry
            word_access_0_1130: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0 
              signal word_access_0_1130_start: Boolean;
              signal Xentry_1131_symbol: Boolean;
              signal Xexit_1132_symbol: Boolean;
              signal cr_1133_symbol : Boolean;
              signal ca_1134_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1130_start <= Xentry_1128_symbol; -- control passed to block
              Xentry_1131_symbol  <= word_access_0_1130_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/$entry
              cr_1133_symbol <= Xentry_1131_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/cr
              simple_obj_ref_289_load_0_req_1 <= cr_1133_symbol; -- link to DP
              ca_1134_symbol <= simple_obj_ref_289_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/ca
              Xexit_1132_symbol <= ca_1134_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0/$exit
              word_access_0_1130_symbol <= Xexit_1132_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/word_access_0
            Xexit_1129_symbol <= word_access_0_1130_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access/$exit
            word_access_1127_symbol <= Xexit_1129_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/word_access
          merge_req_1135_symbol <= word_access_1127_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/merge_req
          simple_obj_ref_289_gather_scatter_req_0 <= merge_req_1135_symbol; -- link to DP
          merge_ack_1136_symbol <= simple_obj_ref_289_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/merge_ack
          Xexit_1126_symbol <= merge_ack_1136_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete/$exit
          simple_obj_ref_289_complete_1124_symbol <= Xexit_1126_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_289_complete
        assign_stmt_297_active_x_x1137_symbol <= binary_296_complete_1149_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_297_active_
        assign_stmt_297_completed_x_x1138_symbol <= assign_stmt_297_active_x_x1137_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/assign_stmt_297_completed_
        binary_296_active_x_x1139_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_active_ 
          signal binary_296_active_x_x1139_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_296_active_x_x1139_predecessors(0) <= binary_296_trigger_x_x1140_symbol;
          binary_296_active_x_x1139_predecessors(1) <= type_cast_293_complete_1144_symbol;
          binary_296_active_x_x1139_join: join -- 
            port map( -- 
              preds => binary_296_active_x_x1139_predecessors,
              symbol_out => binary_296_active_x_x1139_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_active_
        binary_296_trigger_x_x1140_symbol <= Xentry_1043_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_trigger_
        type_cast_293_active_x_x1141_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_active_ 
          signal type_cast_293_active_x_x1141_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_293_active_x_x1141_predecessors(0) <= type_cast_293_trigger_x_x1142_symbol;
          type_cast_293_active_x_x1141_predecessors(1) <= simple_obj_ref_292_complete_1143_symbol;
          type_cast_293_active_x_x1141_join: join -- 
            port map( -- 
              preds => type_cast_293_active_x_x1141_predecessors,
              symbol_out => type_cast_293_active_x_x1141_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_active_
        type_cast_293_trigger_x_x1142_symbol <= Xentry_1043_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_trigger_
        simple_obj_ref_292_complete_1143_symbol <= assign_stmt_290_completed_x_x1108_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/simple_obj_ref_292_complete
        type_cast_293_complete_1144: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete 
          signal type_cast_293_complete_1144_start: Boolean;
          signal Xentry_1145_symbol: Boolean;
          signal Xexit_1146_symbol: Boolean;
          signal req_1147_symbol : Boolean;
          signal ack_1148_symbol : Boolean;
          -- 
        begin -- 
          type_cast_293_complete_1144_start <= type_cast_293_active_x_x1141_symbol; -- control passed to block
          Xentry_1145_symbol  <= type_cast_293_complete_1144_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/$entry
          req_1147_symbol <= Xentry_1145_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/req
          type_cast_293_inst_req_0 <= req_1147_symbol; -- link to DP
          ack_1148_symbol <= type_cast_293_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/ack
          Xexit_1146_symbol <= ack_1148_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete/$exit
          type_cast_293_complete_1144_symbol <= Xexit_1146_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/type_cast_293_complete
        binary_296_complete_1149: Block -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete 
          signal binary_296_complete_1149_start: Boolean;
          signal Xentry_1150_symbol: Boolean;
          signal Xexit_1151_symbol: Boolean;
          signal rr_1152_symbol : Boolean;
          signal ra_1153_symbol : Boolean;
          signal cr_1154_symbol : Boolean;
          signal ca_1155_symbol : Boolean;
          -- 
        begin -- 
          binary_296_complete_1149_start <= binary_296_active_x_x1139_symbol; -- control passed to block
          Xentry_1150_symbol  <= binary_296_complete_1149_start; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/$entry
          rr_1152_symbol <= Xentry_1150_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/rr
          binary_296_inst_req_0 <= rr_1152_symbol; -- link to DP
          ra_1153_symbol <= binary_296_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/ra
          cr_1154_symbol <= ra_1153_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/cr
          binary_296_inst_req_1 <= cr_1154_symbol; -- link to DP
          ca_1155_symbol <= binary_296_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/ca
          Xexit_1151_symbol <= ca_1155_symbol; -- transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete/$exit
          binary_296_complete_1149_symbol <= Xexit_1151_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/binary_296_complete
        Xexit_1044_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/$exit 
          signal Xexit_1044_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          Xexit_1044_predecessors(0) <= assign_stmt_287_completed_x_x1076_symbol;
          Xexit_1044_predecessors(1) <= ptr_deref_285_base_address_calculated_1080_symbol;
          Xexit_1044_predecessors(2) <= assign_stmt_297_completed_x_x1138_symbol;
          Xexit_1044_join: join -- 
            port map( -- 
              preds => Xexit_1044_predecessors,
              symbol_out => Xexit_1044_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297/$exit
        assign_stmt_283_to_assign_stmt_297_1042_symbol <= Xexit_1044_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_283_to_assign_stmt_297
      if_stmt_298_dead_link_1156: Block -- branch_block_stmt_134/if_stmt_298_dead_link 
        signal if_stmt_298_dead_link_1156_start: Boolean;
        signal Xentry_1157_symbol: Boolean;
        signal Xexit_1158_symbol: Boolean;
        signal dead_transition_1159_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_dead_link_1156_start <= if_stmt_298_x_xentry_x_xx_x420_symbol; -- control passed to block
        Xentry_1157_symbol  <= if_stmt_298_dead_link_1156_start; -- transition branch_block_stmt_134/if_stmt_298_dead_link/$entry
        dead_transition_1159_symbol <= false;
        Xexit_1158_symbol <= dead_transition_1159_symbol; -- transition branch_block_stmt_134/if_stmt_298_dead_link/$exit
        if_stmt_298_dead_link_1156_symbol <= Xexit_1158_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_dead_link
      if_stmt_298_eval_test_1160: Block -- branch_block_stmt_134/if_stmt_298_eval_test 
        signal if_stmt_298_eval_test_1160_start: Boolean;
        signal Xentry_1161_symbol: Boolean;
        signal Xexit_1162_symbol: Boolean;
        signal branch_req_1163_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_eval_test_1160_start <= if_stmt_298_x_xentry_x_xx_x420_symbol; -- control passed to block
        Xentry_1161_symbol  <= if_stmt_298_eval_test_1160_start; -- transition branch_block_stmt_134/if_stmt_298_eval_test/$entry
        branch_req_1163_symbol <= Xentry_1161_symbol; -- transition branch_block_stmt_134/if_stmt_298_eval_test/branch_req
        if_stmt_298_branch_req_0 <= branch_req_1163_symbol; -- link to DP
        Xexit_1162_symbol <= branch_req_1163_symbol; -- transition branch_block_stmt_134/if_stmt_298_eval_test/$exit
        if_stmt_298_eval_test_1160_symbol <= Xexit_1162_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_eval_test
      simple_obj_ref_299_place_1164_symbol  <=  if_stmt_298_eval_test_1160_symbol; -- place branch_block_stmt_134/simple_obj_ref_299_place (optimized away) 
      if_stmt_298_if_link_1165: Block -- branch_block_stmt_134/if_stmt_298_if_link 
        signal if_stmt_298_if_link_1165_start: Boolean;
        signal Xentry_1166_symbol: Boolean;
        signal Xexit_1167_symbol: Boolean;
        signal if_choice_transition_1168_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_if_link_1165_start <= simple_obj_ref_299_place_1164_symbol; -- control passed to block
        Xentry_1166_symbol  <= if_stmt_298_if_link_1165_start; -- transition branch_block_stmt_134/if_stmt_298_if_link/$entry
        if_choice_transition_1168_symbol <= if_stmt_298_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_298_if_link/if_choice_transition
        Xexit_1167_symbol <= if_choice_transition_1168_symbol; -- transition branch_block_stmt_134/if_stmt_298_if_link/$exit
        if_stmt_298_if_link_1165_symbol <= Xexit_1167_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_if_link
      if_stmt_298_else_link_1169: Block -- branch_block_stmt_134/if_stmt_298_else_link 
        signal if_stmt_298_else_link_1169_start: Boolean;
        signal Xentry_1170_symbol: Boolean;
        signal Xexit_1171_symbol: Boolean;
        signal else_choice_transition_1172_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_298_else_link_1169_start <= simple_obj_ref_299_place_1164_symbol; -- control passed to block
        Xentry_1170_symbol  <= if_stmt_298_else_link_1169_start; -- transition branch_block_stmt_134/if_stmt_298_else_link/$entry
        else_choice_transition_1172_symbol <= if_stmt_298_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_298_else_link/else_choice_transition
        Xexit_1171_symbol <= else_choice_transition_1172_symbol; -- transition branch_block_stmt_134/if_stmt_298_else_link/$exit
        if_stmt_298_else_link_1169_symbol <= Xexit_1171_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_298_else_link
      bb_5_bb_6_1173_symbol  <=  if_stmt_298_if_link_1165_symbol; -- place branch_block_stmt_134/bb_5_bb_6 (optimized away) 
      bb_5_bb_7_1174_symbol  <=  if_stmt_298_else_link_1169_symbol; -- place branch_block_stmt_134/bb_5_bb_7 (optimized away) 
      assign_stmt_307_to_assign_stmt_319_1175: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319 
        signal assign_stmt_307_to_assign_stmt_319_1175_start: Boolean;
        signal Xentry_1176_symbol: Boolean;
        signal Xexit_1177_symbol: Boolean;
        signal assign_stmt_307_active_x_x1178_symbol : Boolean;
        signal assign_stmt_307_completed_x_x1179_symbol : Boolean;
        signal simple_obj_ref_306_trigger_x_x1180_symbol : Boolean;
        signal simple_obj_ref_306_active_x_x1181_symbol : Boolean;
        signal simple_obj_ref_306_root_address_calculated_1182_symbol : Boolean;
        signal simple_obj_ref_306_word_address_calculated_1183_symbol : Boolean;
        signal simple_obj_ref_306_request_1184_symbol : Boolean;
        signal simple_obj_ref_306_complete_1195_symbol : Boolean;
        signal assign_stmt_312_active_x_x1208_symbol : Boolean;
        signal assign_stmt_312_completed_x_x1209_symbol : Boolean;
        signal array_obj_ref_311_trigger_x_x1210_symbol : Boolean;
        signal array_obj_ref_311_active_x_x1211_symbol : Boolean;
        signal array_obj_ref_311_base_address_calculated_1212_symbol : Boolean;
        signal array_obj_ref_311_root_address_calculated_1213_symbol : Boolean;
        signal array_obj_ref_311_base_address_resized_1214_symbol : Boolean;
        signal array_obj_ref_311_base_addr_resize_1215_symbol : Boolean;
        signal array_obj_ref_311_base_plus_offset_1220_symbol : Boolean;
        signal array_obj_ref_311_complete_1225_symbol : Boolean;
        signal assign_stmt_316_active_x_x1230_symbol : Boolean;
        signal assign_stmt_316_completed_x_x1231_symbol : Boolean;
        signal ptr_deref_315_trigger_x_x1232_symbol : Boolean;
        signal ptr_deref_315_active_x_x1233_symbol : Boolean;
        signal ptr_deref_315_base_address_calculated_1234_symbol : Boolean;
        signal simple_obj_ref_314_complete_1235_symbol : Boolean;
        signal ptr_deref_315_root_address_calculated_1236_symbol : Boolean;
        signal ptr_deref_315_word_address_calculated_1237_symbol : Boolean;
        signal ptr_deref_315_base_address_resized_1238_symbol : Boolean;
        signal ptr_deref_315_base_addr_resize_1239_symbol : Boolean;
        signal ptr_deref_315_base_plus_offset_1244_symbol : Boolean;
        signal ptr_deref_315_word_addrgen_1249_symbol : Boolean;
        signal ptr_deref_315_request_1254_symbol : Boolean;
        signal ptr_deref_315_complete_1265_symbol : Boolean;
        signal assign_stmt_319_active_x_x1278_symbol : Boolean;
        signal assign_stmt_319_completed_x_x1279_symbol : Boolean;
        signal simple_obj_ref_318_complete_1280_symbol : Boolean;
        signal simple_obj_ref_317_trigger_x_x1281_symbol : Boolean;
        signal simple_obj_ref_317_active_x_x1282_symbol : Boolean;
        signal simple_obj_ref_317_root_address_calculated_1283_symbol : Boolean;
        signal simple_obj_ref_317_word_address_calculated_1284_symbol : Boolean;
        signal simple_obj_ref_317_request_1285_symbol : Boolean;
        signal simple_obj_ref_317_complete_1298_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_307_to_assign_stmt_319_1175_start <= assign_stmt_307_to_assign_stmt_319_x_xentry_x_xx_x424_symbol; -- control passed to block
        Xentry_1176_symbol  <= assign_stmt_307_to_assign_stmt_319_1175_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/$entry
        assign_stmt_307_active_x_x1178_symbol <= simple_obj_ref_306_complete_1195_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_307_active_
        assign_stmt_307_completed_x_x1179_symbol <= assign_stmt_307_active_x_x1178_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_307_completed_
        simple_obj_ref_306_trigger_x_x1180_symbol <= simple_obj_ref_306_word_address_calculated_1183_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_trigger_
        simple_obj_ref_306_active_x_x1181_symbol <= simple_obj_ref_306_request_1184_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_active_
        simple_obj_ref_306_root_address_calculated_1182_symbol <= Xentry_1176_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_root_address_calculated
        simple_obj_ref_306_word_address_calculated_1183_symbol <= simple_obj_ref_306_root_address_calculated_1182_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_word_address_calculated
        simple_obj_ref_306_request_1184: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request 
          signal simple_obj_ref_306_request_1184_start: Boolean;
          signal Xentry_1185_symbol: Boolean;
          signal Xexit_1186_symbol: Boolean;
          signal word_access_1187_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_306_request_1184_start <= simple_obj_ref_306_trigger_x_x1180_symbol; -- control passed to block
          Xentry_1185_symbol  <= simple_obj_ref_306_request_1184_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/$entry
          word_access_1187: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access 
            signal word_access_1187_start: Boolean;
            signal Xentry_1188_symbol: Boolean;
            signal Xexit_1189_symbol: Boolean;
            signal word_access_0_1190_symbol : Boolean;
            -- 
          begin -- 
            word_access_1187_start <= Xentry_1185_symbol; -- control passed to block
            Xentry_1188_symbol  <= word_access_1187_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/$entry
            word_access_0_1190: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0 
              signal word_access_0_1190_start: Boolean;
              signal Xentry_1191_symbol: Boolean;
              signal Xexit_1192_symbol: Boolean;
              signal rr_1193_symbol : Boolean;
              signal ra_1194_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1190_start <= Xentry_1188_symbol; -- control passed to block
              Xentry_1191_symbol  <= word_access_0_1190_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/$entry
              rr_1193_symbol <= Xentry_1191_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/rr
              simple_obj_ref_306_load_0_req_0 <= rr_1193_symbol; -- link to DP
              ra_1194_symbol <= simple_obj_ref_306_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/ra
              Xexit_1192_symbol <= ra_1194_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0/$exit
              word_access_0_1190_symbol <= Xexit_1192_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/word_access_0
            Xexit_1189_symbol <= word_access_0_1190_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access/$exit
            word_access_1187_symbol <= Xexit_1189_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/word_access
          Xexit_1186_symbol <= word_access_1187_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request/$exit
          simple_obj_ref_306_request_1184_symbol <= Xexit_1186_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_request
        simple_obj_ref_306_complete_1195: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete 
          signal simple_obj_ref_306_complete_1195_start: Boolean;
          signal Xentry_1196_symbol: Boolean;
          signal Xexit_1197_symbol: Boolean;
          signal word_access_1198_symbol : Boolean;
          signal merge_req_1206_symbol : Boolean;
          signal merge_ack_1207_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_306_complete_1195_start <= simple_obj_ref_306_active_x_x1181_symbol; -- control passed to block
          Xentry_1196_symbol  <= simple_obj_ref_306_complete_1195_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/$entry
          word_access_1198: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access 
            signal word_access_1198_start: Boolean;
            signal Xentry_1199_symbol: Boolean;
            signal Xexit_1200_symbol: Boolean;
            signal word_access_0_1201_symbol : Boolean;
            -- 
          begin -- 
            word_access_1198_start <= Xentry_1196_symbol; -- control passed to block
            Xentry_1199_symbol  <= word_access_1198_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/$entry
            word_access_0_1201: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0 
              signal word_access_0_1201_start: Boolean;
              signal Xentry_1202_symbol: Boolean;
              signal Xexit_1203_symbol: Boolean;
              signal cr_1204_symbol : Boolean;
              signal ca_1205_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1201_start <= Xentry_1199_symbol; -- control passed to block
              Xentry_1202_symbol  <= word_access_0_1201_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/$entry
              cr_1204_symbol <= Xentry_1202_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/cr
              simple_obj_ref_306_load_0_req_1 <= cr_1204_symbol; -- link to DP
              ca_1205_symbol <= simple_obj_ref_306_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/ca
              Xexit_1203_symbol <= ca_1205_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0/$exit
              word_access_0_1201_symbol <= Xexit_1203_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/word_access_0
            Xexit_1200_symbol <= word_access_0_1201_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access/$exit
            word_access_1198_symbol <= Xexit_1200_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/word_access
          merge_req_1206_symbol <= word_access_1198_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/merge_req
          simple_obj_ref_306_gather_scatter_req_0 <= merge_req_1206_symbol; -- link to DP
          merge_ack_1207_symbol <= simple_obj_ref_306_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/merge_ack
          Xexit_1197_symbol <= merge_ack_1207_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete/$exit
          simple_obj_ref_306_complete_1195_symbol <= Xexit_1197_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_306_complete
        assign_stmt_312_active_x_x1208_symbol <= array_obj_ref_311_complete_1225_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_312_active_
        assign_stmt_312_completed_x_x1209_symbol <= assign_stmt_312_active_x_x1208_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_312_completed_
        array_obj_ref_311_trigger_x_x1210_symbol <= Xentry_1176_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_trigger_
        array_obj_ref_311_active_x_x1211_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_active_ 
          signal array_obj_ref_311_active_x_x1211_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_311_active_x_x1211_predecessors(0) <= array_obj_ref_311_trigger_x_x1210_symbol;
          array_obj_ref_311_active_x_x1211_predecessors(1) <= array_obj_ref_311_root_address_calculated_1213_symbol;
          array_obj_ref_311_active_x_x1211_join: join -- 
            port map( -- 
              preds => array_obj_ref_311_active_x_x1211_predecessors,
              symbol_out => array_obj_ref_311_active_x_x1211_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_active_
        array_obj_ref_311_base_address_calculated_1212_symbol <= assign_stmt_307_completed_x_x1179_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_address_calculated
        array_obj_ref_311_root_address_calculated_1213_symbol <= array_obj_ref_311_base_plus_offset_1220_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_root_address_calculated
        array_obj_ref_311_base_address_resized_1214_symbol <= array_obj_ref_311_base_addr_resize_1215_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_address_resized
        array_obj_ref_311_base_addr_resize_1215: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize 
          signal array_obj_ref_311_base_addr_resize_1215_start: Boolean;
          signal Xentry_1216_symbol: Boolean;
          signal Xexit_1217_symbol: Boolean;
          signal base_resize_req_1218_symbol : Boolean;
          signal base_resize_ack_1219_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_311_base_addr_resize_1215_start <= array_obj_ref_311_base_address_calculated_1212_symbol; -- control passed to block
          Xentry_1216_symbol  <= array_obj_ref_311_base_addr_resize_1215_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/$entry
          base_resize_req_1218_symbol <= Xentry_1216_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/base_resize_req
          array_obj_ref_311_base_resize_req_0 <= base_resize_req_1218_symbol; -- link to DP
          base_resize_ack_1219_symbol <= array_obj_ref_311_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/base_resize_ack
          Xexit_1217_symbol <= base_resize_ack_1219_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize/$exit
          array_obj_ref_311_base_addr_resize_1215_symbol <= Xexit_1217_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_addr_resize
        array_obj_ref_311_base_plus_offset_1220: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset 
          signal array_obj_ref_311_base_plus_offset_1220_start: Boolean;
          signal Xentry_1221_symbol: Boolean;
          signal Xexit_1222_symbol: Boolean;
          signal sum_rename_req_1223_symbol : Boolean;
          signal sum_rename_ack_1224_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_311_base_plus_offset_1220_start <= array_obj_ref_311_base_address_resized_1214_symbol; -- control passed to block
          Xentry_1221_symbol  <= array_obj_ref_311_base_plus_offset_1220_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/$entry
          sum_rename_req_1223_symbol <= Xentry_1221_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/sum_rename_req
          array_obj_ref_311_root_address_inst_req_0 <= sum_rename_req_1223_symbol; -- link to DP
          sum_rename_ack_1224_symbol <= array_obj_ref_311_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/sum_rename_ack
          Xexit_1222_symbol <= sum_rename_ack_1224_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset/$exit
          array_obj_ref_311_base_plus_offset_1220_symbol <= Xexit_1222_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_base_plus_offset
        array_obj_ref_311_complete_1225: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete 
          signal array_obj_ref_311_complete_1225_start: Boolean;
          signal Xentry_1226_symbol: Boolean;
          signal Xexit_1227_symbol: Boolean;
          signal final_reg_req_1228_symbol : Boolean;
          signal final_reg_ack_1229_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_311_complete_1225_start <= array_obj_ref_311_active_x_x1211_symbol; -- control passed to block
          Xentry_1226_symbol  <= array_obj_ref_311_complete_1225_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/$entry
          final_reg_req_1228_symbol <= Xentry_1226_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/final_reg_req
          array_obj_ref_311_final_reg_req_0 <= final_reg_req_1228_symbol; -- link to DP
          final_reg_ack_1229_symbol <= array_obj_ref_311_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/final_reg_ack
          Xexit_1227_symbol <= final_reg_ack_1229_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete/$exit
          array_obj_ref_311_complete_1225_symbol <= Xexit_1227_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/array_obj_ref_311_complete
        assign_stmt_316_active_x_x1230_symbol <= ptr_deref_315_complete_1265_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_316_active_
        assign_stmt_316_completed_x_x1231_symbol <= assign_stmt_316_active_x_x1230_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_316_completed_
        ptr_deref_315_trigger_x_x1232_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_trigger_ 
          signal ptr_deref_315_trigger_x_x1232_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_315_trigger_x_x1232_predecessors(0) <= ptr_deref_315_word_address_calculated_1237_symbol;
          ptr_deref_315_trigger_x_x1232_predecessors(1) <= ptr_deref_315_base_address_calculated_1234_symbol;
          ptr_deref_315_trigger_x_x1232_join: join -- 
            port map( -- 
              preds => ptr_deref_315_trigger_x_x1232_predecessors,
              symbol_out => ptr_deref_315_trigger_x_x1232_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_trigger_
        ptr_deref_315_active_x_x1233_symbol <= ptr_deref_315_request_1254_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_active_
        ptr_deref_315_base_address_calculated_1234_symbol <= simple_obj_ref_314_complete_1235_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_address_calculated
        simple_obj_ref_314_complete_1235_symbol <= assign_stmt_312_completed_x_x1209_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_314_complete
        ptr_deref_315_root_address_calculated_1236_symbol <= ptr_deref_315_base_plus_offset_1244_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_root_address_calculated
        ptr_deref_315_word_address_calculated_1237_symbol <= ptr_deref_315_word_addrgen_1249_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_address_calculated
        ptr_deref_315_base_address_resized_1238_symbol <= ptr_deref_315_base_addr_resize_1239_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_address_resized
        ptr_deref_315_base_addr_resize_1239: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize 
          signal ptr_deref_315_base_addr_resize_1239_start: Boolean;
          signal Xentry_1240_symbol: Boolean;
          signal Xexit_1241_symbol: Boolean;
          signal base_resize_req_1242_symbol : Boolean;
          signal base_resize_ack_1243_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_base_addr_resize_1239_start <= ptr_deref_315_base_address_calculated_1234_symbol; -- control passed to block
          Xentry_1240_symbol  <= ptr_deref_315_base_addr_resize_1239_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/$entry
          base_resize_req_1242_symbol <= Xentry_1240_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/base_resize_req
          ptr_deref_315_base_resize_req_0 <= base_resize_req_1242_symbol; -- link to DP
          base_resize_ack_1243_symbol <= ptr_deref_315_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/base_resize_ack
          Xexit_1241_symbol <= base_resize_ack_1243_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize/$exit
          ptr_deref_315_base_addr_resize_1239_symbol <= Xexit_1241_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_addr_resize
        ptr_deref_315_base_plus_offset_1244: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset 
          signal ptr_deref_315_base_plus_offset_1244_start: Boolean;
          signal Xentry_1245_symbol: Boolean;
          signal Xexit_1246_symbol: Boolean;
          signal sum_rename_req_1247_symbol : Boolean;
          signal sum_rename_ack_1248_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_base_plus_offset_1244_start <= ptr_deref_315_base_address_resized_1238_symbol; -- control passed to block
          Xentry_1245_symbol  <= ptr_deref_315_base_plus_offset_1244_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/$entry
          sum_rename_req_1247_symbol <= Xentry_1245_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/sum_rename_req
          ptr_deref_315_root_address_inst_req_0 <= sum_rename_req_1247_symbol; -- link to DP
          sum_rename_ack_1248_symbol <= ptr_deref_315_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/sum_rename_ack
          Xexit_1246_symbol <= sum_rename_ack_1248_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset/$exit
          ptr_deref_315_base_plus_offset_1244_symbol <= Xexit_1246_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_base_plus_offset
        ptr_deref_315_word_addrgen_1249: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen 
          signal ptr_deref_315_word_addrgen_1249_start: Boolean;
          signal Xentry_1250_symbol: Boolean;
          signal Xexit_1251_symbol: Boolean;
          signal root_rename_req_1252_symbol : Boolean;
          signal root_rename_ack_1253_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_word_addrgen_1249_start <= ptr_deref_315_root_address_calculated_1236_symbol; -- control passed to block
          Xentry_1250_symbol  <= ptr_deref_315_word_addrgen_1249_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/$entry
          root_rename_req_1252_symbol <= Xentry_1250_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/root_rename_req
          ptr_deref_315_addr_0_req_0 <= root_rename_req_1252_symbol; -- link to DP
          root_rename_ack_1253_symbol <= ptr_deref_315_addr_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/root_rename_ack
          Xexit_1251_symbol <= root_rename_ack_1253_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen/$exit
          ptr_deref_315_word_addrgen_1249_symbol <= Xexit_1251_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_word_addrgen
        ptr_deref_315_request_1254: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request 
          signal ptr_deref_315_request_1254_start: Boolean;
          signal Xentry_1255_symbol: Boolean;
          signal Xexit_1256_symbol: Boolean;
          signal word_access_1257_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_request_1254_start <= ptr_deref_315_trigger_x_x1232_symbol; -- control passed to block
          Xentry_1255_symbol  <= ptr_deref_315_request_1254_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/$entry
          word_access_1257: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access 
            signal word_access_1257_start: Boolean;
            signal Xentry_1258_symbol: Boolean;
            signal Xexit_1259_symbol: Boolean;
            signal word_access_0_1260_symbol : Boolean;
            -- 
          begin -- 
            word_access_1257_start <= Xentry_1255_symbol; -- control passed to block
            Xentry_1258_symbol  <= word_access_1257_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/$entry
            word_access_0_1260: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0 
              signal word_access_0_1260_start: Boolean;
              signal Xentry_1261_symbol: Boolean;
              signal Xexit_1262_symbol: Boolean;
              signal rr_1263_symbol : Boolean;
              signal ra_1264_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1260_start <= Xentry_1258_symbol; -- control passed to block
              Xentry_1261_symbol  <= word_access_0_1260_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/$entry
              rr_1263_symbol <= Xentry_1261_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/rr
              ptr_deref_315_load_0_req_0 <= rr_1263_symbol; -- link to DP
              ra_1264_symbol <= ptr_deref_315_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/ra
              Xexit_1262_symbol <= ra_1264_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0/$exit
              word_access_0_1260_symbol <= Xexit_1262_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/word_access_0
            Xexit_1259_symbol <= word_access_0_1260_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access/$exit
            word_access_1257_symbol <= Xexit_1259_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/word_access
          Xexit_1256_symbol <= word_access_1257_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request/$exit
          ptr_deref_315_request_1254_symbol <= Xexit_1256_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_request
        ptr_deref_315_complete_1265: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete 
          signal ptr_deref_315_complete_1265_start: Boolean;
          signal Xentry_1266_symbol: Boolean;
          signal Xexit_1267_symbol: Boolean;
          signal word_access_1268_symbol : Boolean;
          signal merge_req_1276_symbol : Boolean;
          signal merge_ack_1277_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_315_complete_1265_start <= ptr_deref_315_active_x_x1233_symbol; -- control passed to block
          Xentry_1266_symbol  <= ptr_deref_315_complete_1265_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/$entry
          word_access_1268: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access 
            signal word_access_1268_start: Boolean;
            signal Xentry_1269_symbol: Boolean;
            signal Xexit_1270_symbol: Boolean;
            signal word_access_0_1271_symbol : Boolean;
            -- 
          begin -- 
            word_access_1268_start <= Xentry_1266_symbol; -- control passed to block
            Xentry_1269_symbol  <= word_access_1268_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/$entry
            word_access_0_1271: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0 
              signal word_access_0_1271_start: Boolean;
              signal Xentry_1272_symbol: Boolean;
              signal Xexit_1273_symbol: Boolean;
              signal cr_1274_symbol : Boolean;
              signal ca_1275_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1271_start <= Xentry_1269_symbol; -- control passed to block
              Xentry_1272_symbol  <= word_access_0_1271_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/$entry
              cr_1274_symbol <= Xentry_1272_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/cr
              ptr_deref_315_load_0_req_1 <= cr_1274_symbol; -- link to DP
              ca_1275_symbol <= ptr_deref_315_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/ca
              Xexit_1273_symbol <= ca_1275_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0/$exit
              word_access_0_1271_symbol <= Xexit_1273_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/word_access_0
            Xexit_1270_symbol <= word_access_0_1271_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access/$exit
            word_access_1268_symbol <= Xexit_1270_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/word_access
          merge_req_1276_symbol <= word_access_1268_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/merge_req
          ptr_deref_315_gather_scatter_req_0 <= merge_req_1276_symbol; -- link to DP
          merge_ack_1277_symbol <= ptr_deref_315_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/merge_ack
          Xexit_1267_symbol <= merge_ack_1277_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete/$exit
          ptr_deref_315_complete_1265_symbol <= Xexit_1267_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/ptr_deref_315_complete
        assign_stmt_319_active_x_x1278_symbol <= simple_obj_ref_318_complete_1280_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_319_active_
        assign_stmt_319_completed_x_x1279_symbol <= simple_obj_ref_317_complete_1298_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/assign_stmt_319_completed_
        simple_obj_ref_318_complete_1280_symbol <= assign_stmt_316_completed_x_x1231_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_318_complete
        simple_obj_ref_317_trigger_x_x1281_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_trigger_ 
          signal simple_obj_ref_317_trigger_x_x1281_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          simple_obj_ref_317_trigger_x_x1281_predecessors(0) <= simple_obj_ref_317_word_address_calculated_1284_symbol;
          simple_obj_ref_317_trigger_x_x1281_predecessors(1) <= assign_stmt_319_active_x_x1278_symbol;
          simple_obj_ref_317_trigger_x_x1281_predecessors(2) <= simple_obj_ref_306_active_x_x1181_symbol;
          simple_obj_ref_317_trigger_x_x1281_join: join -- 
            port map( -- 
              preds => simple_obj_ref_317_trigger_x_x1281_predecessors,
              symbol_out => simple_obj_ref_317_trigger_x_x1281_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_trigger_
        simple_obj_ref_317_active_x_x1282_symbol <= simple_obj_ref_317_request_1285_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_active_
        simple_obj_ref_317_root_address_calculated_1283_symbol <= Xentry_1176_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_root_address_calculated
        simple_obj_ref_317_word_address_calculated_1284_symbol <= simple_obj_ref_317_root_address_calculated_1283_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_word_address_calculated
        simple_obj_ref_317_request_1285: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request 
          signal simple_obj_ref_317_request_1285_start: Boolean;
          signal Xentry_1286_symbol: Boolean;
          signal Xexit_1287_symbol: Boolean;
          signal split_req_1288_symbol : Boolean;
          signal split_ack_1289_symbol : Boolean;
          signal word_access_1290_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_317_request_1285_start <= simple_obj_ref_317_trigger_x_x1281_symbol; -- control passed to block
          Xentry_1286_symbol  <= simple_obj_ref_317_request_1285_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/$entry
          split_req_1288_symbol <= Xentry_1286_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/split_req
          simple_obj_ref_317_gather_scatter_req_0 <= split_req_1288_symbol; -- link to DP
          split_ack_1289_symbol <= simple_obj_ref_317_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/split_ack
          word_access_1290: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access 
            signal word_access_1290_start: Boolean;
            signal Xentry_1291_symbol: Boolean;
            signal Xexit_1292_symbol: Boolean;
            signal word_access_0_1293_symbol : Boolean;
            -- 
          begin -- 
            word_access_1290_start <= split_ack_1289_symbol; -- control passed to block
            Xentry_1291_symbol  <= word_access_1290_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/$entry
            word_access_0_1293: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0 
              signal word_access_0_1293_start: Boolean;
              signal Xentry_1294_symbol: Boolean;
              signal Xexit_1295_symbol: Boolean;
              signal rr_1296_symbol : Boolean;
              signal ra_1297_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1293_start <= Xentry_1291_symbol; -- control passed to block
              Xentry_1294_symbol  <= word_access_0_1293_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/$entry
              rr_1296_symbol <= Xentry_1294_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/rr
              simple_obj_ref_317_store_0_req_0 <= rr_1296_symbol; -- link to DP
              ra_1297_symbol <= simple_obj_ref_317_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/ra
              Xexit_1295_symbol <= ra_1297_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0/$exit
              word_access_0_1293_symbol <= Xexit_1295_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/word_access_0
            Xexit_1292_symbol <= word_access_0_1293_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access/$exit
            word_access_1290_symbol <= Xexit_1292_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/word_access
          Xexit_1287_symbol <= word_access_1290_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request/$exit
          simple_obj_ref_317_request_1285_symbol <= Xexit_1287_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_request
        simple_obj_ref_317_complete_1298: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete 
          signal simple_obj_ref_317_complete_1298_start: Boolean;
          signal Xentry_1299_symbol: Boolean;
          signal Xexit_1300_symbol: Boolean;
          signal word_access_1301_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_317_complete_1298_start <= simple_obj_ref_317_active_x_x1282_symbol; -- control passed to block
          Xentry_1299_symbol  <= simple_obj_ref_317_complete_1298_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/$entry
          word_access_1301: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access 
            signal word_access_1301_start: Boolean;
            signal Xentry_1302_symbol: Boolean;
            signal Xexit_1303_symbol: Boolean;
            signal word_access_0_1304_symbol : Boolean;
            -- 
          begin -- 
            word_access_1301_start <= Xentry_1299_symbol; -- control passed to block
            Xentry_1302_symbol  <= word_access_1301_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/$entry
            word_access_0_1304: Block -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0 
              signal word_access_0_1304_start: Boolean;
              signal Xentry_1305_symbol: Boolean;
              signal Xexit_1306_symbol: Boolean;
              signal cr_1307_symbol : Boolean;
              signal ca_1308_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1304_start <= Xentry_1302_symbol; -- control passed to block
              Xentry_1305_symbol  <= word_access_0_1304_start; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/$entry
              cr_1307_symbol <= Xentry_1305_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/cr
              simple_obj_ref_317_store_0_req_1 <= cr_1307_symbol; -- link to DP
              ca_1308_symbol <= simple_obj_ref_317_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/ca
              Xexit_1306_symbol <= ca_1308_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0/$exit
              word_access_0_1304_symbol <= Xexit_1306_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/word_access_0
            Xexit_1303_symbol <= word_access_0_1304_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access/$exit
            word_access_1301_symbol <= Xexit_1303_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/word_access
          Xexit_1300_symbol <= word_access_1301_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete/$exit
          simple_obj_ref_317_complete_1298_symbol <= Xexit_1300_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/simple_obj_ref_317_complete
        Xexit_1177_symbol <= assign_stmt_319_completed_x_x1279_symbol; -- transition branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319/$exit
        assign_stmt_307_to_assign_stmt_319_1175_symbol <= Xexit_1177_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_307_to_assign_stmt_319
      assign_stmt_325_to_assign_stmt_334_1309: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334 
        signal assign_stmt_325_to_assign_stmt_334_1309_start: Boolean;
        signal Xentry_1310_symbol: Boolean;
        signal Xexit_1311_symbol: Boolean;
        signal assign_stmt_325_active_x_x1312_symbol : Boolean;
        signal assign_stmt_325_completed_x_x1313_symbol : Boolean;
        signal ptr_deref_324_trigger_x_x1314_symbol : Boolean;
        signal ptr_deref_324_active_x_x1315_symbol : Boolean;
        signal ptr_deref_324_base_address_calculated_1316_symbol : Boolean;
        signal ptr_deref_324_root_address_calculated_1317_symbol : Boolean;
        signal ptr_deref_324_word_address_calculated_1318_symbol : Boolean;
        signal ptr_deref_324_request_1319_symbol : Boolean;
        signal ptr_deref_324_complete_1330_symbol : Boolean;
        signal assign_stmt_329_active_x_x1343_symbol : Boolean;
        signal assign_stmt_329_completed_x_x1344_symbol : Boolean;
        signal type_cast_328_active_x_x1345_symbol : Boolean;
        signal type_cast_328_trigger_x_x1346_symbol : Boolean;
        signal simple_obj_ref_327_complete_1347_symbol : Boolean;
        signal type_cast_328_complete_1348_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_325_to_assign_stmt_334_1309_start <= assign_stmt_325_to_assign_stmt_334_x_xentry_x_xx_x428_symbol; -- control passed to block
        Xentry_1310_symbol  <= assign_stmt_325_to_assign_stmt_334_1309_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/$entry
        assign_stmt_325_active_x_x1312_symbol <= ptr_deref_324_complete_1330_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_325_active_
        assign_stmt_325_completed_x_x1313_symbol <= assign_stmt_325_active_x_x1312_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_325_completed_
        ptr_deref_324_trigger_x_x1314_symbol <= ptr_deref_324_word_address_calculated_1318_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_trigger_
        ptr_deref_324_active_x_x1315_symbol <= ptr_deref_324_request_1319_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_active_
        ptr_deref_324_base_address_calculated_1316_symbol <= Xentry_1310_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_base_address_calculated
        ptr_deref_324_root_address_calculated_1317_symbol <= Xentry_1310_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_root_address_calculated
        ptr_deref_324_word_address_calculated_1318_symbol <= ptr_deref_324_root_address_calculated_1317_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_word_address_calculated
        ptr_deref_324_request_1319: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request 
          signal ptr_deref_324_request_1319_start: Boolean;
          signal Xentry_1320_symbol: Boolean;
          signal Xexit_1321_symbol: Boolean;
          signal word_access_1322_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_324_request_1319_start <= ptr_deref_324_trigger_x_x1314_symbol; -- control passed to block
          Xentry_1320_symbol  <= ptr_deref_324_request_1319_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/$entry
          word_access_1322: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access 
            signal word_access_1322_start: Boolean;
            signal Xentry_1323_symbol: Boolean;
            signal Xexit_1324_symbol: Boolean;
            signal word_access_0_1325_symbol : Boolean;
            -- 
          begin -- 
            word_access_1322_start <= Xentry_1320_symbol; -- control passed to block
            Xentry_1323_symbol  <= word_access_1322_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/$entry
            word_access_0_1325: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0 
              signal word_access_0_1325_start: Boolean;
              signal Xentry_1326_symbol: Boolean;
              signal Xexit_1327_symbol: Boolean;
              signal rr_1328_symbol : Boolean;
              signal ra_1329_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1325_start <= Xentry_1323_symbol; -- control passed to block
              Xentry_1326_symbol  <= word_access_0_1325_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/$entry
              rr_1328_symbol <= Xentry_1326_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/rr
              ptr_deref_324_load_0_req_0 <= rr_1328_symbol; -- link to DP
              ra_1329_symbol <= ptr_deref_324_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/ra
              Xexit_1327_symbol <= ra_1329_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0/$exit
              word_access_0_1325_symbol <= Xexit_1327_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/word_access_0
            Xexit_1324_symbol <= word_access_0_1325_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access/$exit
            word_access_1322_symbol <= Xexit_1324_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/word_access
          Xexit_1321_symbol <= word_access_1322_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request/$exit
          ptr_deref_324_request_1319_symbol <= Xexit_1321_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_request
        ptr_deref_324_complete_1330: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete 
          signal ptr_deref_324_complete_1330_start: Boolean;
          signal Xentry_1331_symbol: Boolean;
          signal Xexit_1332_symbol: Boolean;
          signal word_access_1333_symbol : Boolean;
          signal merge_req_1341_symbol : Boolean;
          signal merge_ack_1342_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_324_complete_1330_start <= ptr_deref_324_active_x_x1315_symbol; -- control passed to block
          Xentry_1331_symbol  <= ptr_deref_324_complete_1330_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/$entry
          word_access_1333: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access 
            signal word_access_1333_start: Boolean;
            signal Xentry_1334_symbol: Boolean;
            signal Xexit_1335_symbol: Boolean;
            signal word_access_0_1336_symbol : Boolean;
            -- 
          begin -- 
            word_access_1333_start <= Xentry_1331_symbol; -- control passed to block
            Xentry_1334_symbol  <= word_access_1333_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/$entry
            word_access_0_1336: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0 
              signal word_access_0_1336_start: Boolean;
              signal Xentry_1337_symbol: Boolean;
              signal Xexit_1338_symbol: Boolean;
              signal cr_1339_symbol : Boolean;
              signal ca_1340_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1336_start <= Xentry_1334_symbol; -- control passed to block
              Xentry_1337_symbol  <= word_access_0_1336_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/$entry
              cr_1339_symbol <= Xentry_1337_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/cr
              ptr_deref_324_load_0_req_1 <= cr_1339_symbol; -- link to DP
              ca_1340_symbol <= ptr_deref_324_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/ca
              Xexit_1338_symbol <= ca_1340_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0/$exit
              word_access_0_1336_symbol <= Xexit_1338_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/word_access_0
            Xexit_1335_symbol <= word_access_0_1336_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access/$exit
            word_access_1333_symbol <= Xexit_1335_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/word_access
          merge_req_1341_symbol <= word_access_1333_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/merge_req
          ptr_deref_324_gather_scatter_req_0 <= merge_req_1341_symbol; -- link to DP
          merge_ack_1342_symbol <= ptr_deref_324_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/merge_ack
          Xexit_1332_symbol <= merge_ack_1342_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete/$exit
          ptr_deref_324_complete_1330_symbol <= Xexit_1332_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/ptr_deref_324_complete
        assign_stmt_329_active_x_x1343_symbol <= type_cast_328_complete_1348_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_329_active_
        assign_stmt_329_completed_x_x1344_symbol <= assign_stmt_329_active_x_x1343_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/assign_stmt_329_completed_
        type_cast_328_active_x_x1345_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_active_ 
          signal type_cast_328_active_x_x1345_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_328_active_x_x1345_predecessors(0) <= type_cast_328_trigger_x_x1346_symbol;
          type_cast_328_active_x_x1345_predecessors(1) <= simple_obj_ref_327_complete_1347_symbol;
          type_cast_328_active_x_x1345_join: join -- 
            port map( -- 
              preds => type_cast_328_active_x_x1345_predecessors,
              symbol_out => type_cast_328_active_x_x1345_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_active_
        type_cast_328_trigger_x_x1346_symbol <= Xentry_1310_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_trigger_
        simple_obj_ref_327_complete_1347_symbol <= assign_stmt_325_completed_x_x1313_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/simple_obj_ref_327_complete
        type_cast_328_complete_1348: Block -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete 
          signal type_cast_328_complete_1348_start: Boolean;
          signal Xentry_1349_symbol: Boolean;
          signal Xexit_1350_symbol: Boolean;
          signal req_1351_symbol : Boolean;
          signal ack_1352_symbol : Boolean;
          -- 
        begin -- 
          type_cast_328_complete_1348_start <= type_cast_328_active_x_x1345_symbol; -- control passed to block
          Xentry_1349_symbol  <= type_cast_328_complete_1348_start; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/$entry
          req_1351_symbol <= Xentry_1349_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/req
          type_cast_328_inst_req_0 <= req_1351_symbol; -- link to DP
          ack_1352_symbol <= type_cast_328_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/ack
          Xexit_1350_symbol <= ack_1352_symbol; -- transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete/$exit
          type_cast_328_complete_1348_symbol <= Xexit_1350_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/type_cast_328_complete
        Xexit_1311_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/$exit 
          signal Xexit_1311_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_1311_predecessors(0) <= ptr_deref_324_base_address_calculated_1316_symbol;
          Xexit_1311_predecessors(1) <= assign_stmt_329_completed_x_x1344_symbol;
          Xexit_1311_join: join -- 
            port map( -- 
              preds => Xexit_1311_predecessors,
              symbol_out => Xexit_1311_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334/$exit
        assign_stmt_325_to_assign_stmt_334_1309_symbol <= Xexit_1311_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_325_to_assign_stmt_334
      assign_stmt_338_1353: Block -- branch_block_stmt_134/assign_stmt_338 
        signal assign_stmt_338_1353_start: Boolean;
        signal Xentry_1354_symbol: Boolean;
        signal Xexit_1355_symbol: Boolean;
        signal assign_stmt_338_active_x_x1356_symbol : Boolean;
        signal assign_stmt_338_completed_x_x1357_symbol : Boolean;
        signal type_cast_337_active_x_x1358_symbol : Boolean;
        signal type_cast_337_trigger_x_x1359_symbol : Boolean;
        signal simple_obj_ref_336_complete_1360_symbol : Boolean;
        signal type_cast_337_complete_1361_symbol : Boolean;
        signal simple_obj_ref_335_trigger_x_x1366_symbol : Boolean;
        signal simple_obj_ref_335_complete_1367_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_338_1353_start <= assign_stmt_338_x_xentry_x_xx_x430_symbol; -- control passed to block
        Xentry_1354_symbol  <= assign_stmt_338_1353_start; -- transition branch_block_stmt_134/assign_stmt_338/$entry
        assign_stmt_338_active_x_x1356_symbol <= type_cast_337_complete_1361_symbol; -- transition branch_block_stmt_134/assign_stmt_338/assign_stmt_338_active_
        assign_stmt_338_completed_x_x1357_symbol <= simple_obj_ref_335_complete_1367_symbol; -- transition branch_block_stmt_134/assign_stmt_338/assign_stmt_338_completed_
        type_cast_337_active_x_x1358_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_338/type_cast_337_active_ 
          signal type_cast_337_active_x_x1358_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_337_active_x_x1358_predecessors(0) <= type_cast_337_trigger_x_x1359_symbol;
          type_cast_337_active_x_x1358_predecessors(1) <= simple_obj_ref_336_complete_1360_symbol;
          type_cast_337_active_x_x1358_join: join -- 
            port map( -- 
              preds => type_cast_337_active_x_x1358_predecessors,
              symbol_out => type_cast_337_active_x_x1358_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_338/type_cast_337_active_
        type_cast_337_trigger_x_x1359_symbol <= Xentry_1354_symbol; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_trigger_
        simple_obj_ref_336_complete_1360_symbol <= Xentry_1354_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_336_complete
        type_cast_337_complete_1361: Block -- branch_block_stmt_134/assign_stmt_338/type_cast_337_complete 
          signal type_cast_337_complete_1361_start: Boolean;
          signal Xentry_1362_symbol: Boolean;
          signal Xexit_1363_symbol: Boolean;
          signal req_1364_symbol : Boolean;
          signal ack_1365_symbol : Boolean;
          -- 
        begin -- 
          type_cast_337_complete_1361_start <= type_cast_337_active_x_x1358_symbol; -- control passed to block
          Xentry_1362_symbol  <= type_cast_337_complete_1361_start; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/$entry
          req_1364_symbol <= Xentry_1362_symbol; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/req
          type_cast_337_inst_req_0 <= req_1364_symbol; -- link to DP
          ack_1365_symbol <= type_cast_337_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/ack
          Xexit_1363_symbol <= ack_1365_symbol; -- transition branch_block_stmt_134/assign_stmt_338/type_cast_337_complete/$exit
          type_cast_337_complete_1361_symbol <= Xexit_1363_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_338/type_cast_337_complete
        simple_obj_ref_335_trigger_x_x1366_symbol <= assign_stmt_338_active_x_x1356_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_trigger_
        simple_obj_ref_335_complete_1367: Block -- branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete 
          signal simple_obj_ref_335_complete_1367_start: Boolean;
          signal Xentry_1368_symbol: Boolean;
          signal Xexit_1369_symbol: Boolean;
          signal pipe_wreq_1370_symbol : Boolean;
          signal pipe_wack_1371_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_335_complete_1367_start <= simple_obj_ref_335_trigger_x_x1366_symbol; -- control passed to block
          Xentry_1368_symbol  <= simple_obj_ref_335_complete_1367_start; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/$entry
          pipe_wreq_1370_symbol <= Xentry_1368_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/pipe_wreq
          simple_obj_ref_335_inst_req_0 <= pipe_wreq_1370_symbol; -- link to DP
          pipe_wack_1371_symbol <= simple_obj_ref_335_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/pipe_wack
          Xexit_1369_symbol <= pipe_wack_1371_symbol; -- transition branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete/$exit
          simple_obj_ref_335_complete_1367_symbol <= Xexit_1369_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_338/simple_obj_ref_335_complete
        Xexit_1355_symbol <= assign_stmt_338_completed_x_x1357_symbol; -- transition branch_block_stmt_134/assign_stmt_338/$exit
        assign_stmt_338_1353_symbol <= Xexit_1355_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_338
      assign_stmt_344_to_assign_stmt_353_1372: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353 
        signal assign_stmt_344_to_assign_stmt_353_1372_start: Boolean;
        signal Xentry_1373_symbol: Boolean;
        signal Xexit_1374_symbol: Boolean;
        signal assign_stmt_344_active_x_x1375_symbol : Boolean;
        signal assign_stmt_344_completed_x_x1376_symbol : Boolean;
        signal ptr_deref_343_trigger_x_x1377_symbol : Boolean;
        signal ptr_deref_343_active_x_x1378_symbol : Boolean;
        signal ptr_deref_343_base_address_calculated_1379_symbol : Boolean;
        signal ptr_deref_343_root_address_calculated_1380_symbol : Boolean;
        signal ptr_deref_343_word_address_calculated_1381_symbol : Boolean;
        signal ptr_deref_343_request_1382_symbol : Boolean;
        signal ptr_deref_343_complete_1393_symbol : Boolean;
        signal assign_stmt_348_active_x_x1406_symbol : Boolean;
        signal assign_stmt_348_completed_x_x1407_symbol : Boolean;
        signal type_cast_347_active_x_x1408_symbol : Boolean;
        signal type_cast_347_trigger_x_x1409_symbol : Boolean;
        signal simple_obj_ref_346_complete_1410_symbol : Boolean;
        signal type_cast_347_complete_1411_symbol : Boolean;
        signal assign_stmt_353_active_x_x1416_symbol : Boolean;
        signal assign_stmt_353_completed_x_x1417_symbol : Boolean;
        signal binary_352_active_x_x1418_symbol : Boolean;
        signal binary_352_trigger_x_x1419_symbol : Boolean;
        signal simple_obj_ref_350_complete_1420_symbol : Boolean;
        signal binary_352_complete_1421_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_344_to_assign_stmt_353_1372_start <= assign_stmt_344_to_assign_stmt_353_x_xentry_x_xx_x434_symbol; -- control passed to block
        Xentry_1373_symbol  <= assign_stmt_344_to_assign_stmt_353_1372_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/$entry
        assign_stmt_344_active_x_x1375_symbol <= ptr_deref_343_complete_1393_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_344_active_
        assign_stmt_344_completed_x_x1376_symbol <= assign_stmt_344_active_x_x1375_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_344_completed_
        ptr_deref_343_trigger_x_x1377_symbol <= ptr_deref_343_word_address_calculated_1381_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_trigger_
        ptr_deref_343_active_x_x1378_symbol <= ptr_deref_343_request_1382_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_active_
        ptr_deref_343_base_address_calculated_1379_symbol <= Xentry_1373_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_base_address_calculated
        ptr_deref_343_root_address_calculated_1380_symbol <= Xentry_1373_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_root_address_calculated
        ptr_deref_343_word_address_calculated_1381_symbol <= ptr_deref_343_root_address_calculated_1380_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_word_address_calculated
        ptr_deref_343_request_1382: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request 
          signal ptr_deref_343_request_1382_start: Boolean;
          signal Xentry_1383_symbol: Boolean;
          signal Xexit_1384_symbol: Boolean;
          signal word_access_1385_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_343_request_1382_start <= ptr_deref_343_trigger_x_x1377_symbol; -- control passed to block
          Xentry_1383_symbol  <= ptr_deref_343_request_1382_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/$entry
          word_access_1385: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access 
            signal word_access_1385_start: Boolean;
            signal Xentry_1386_symbol: Boolean;
            signal Xexit_1387_symbol: Boolean;
            signal word_access_0_1388_symbol : Boolean;
            -- 
          begin -- 
            word_access_1385_start <= Xentry_1383_symbol; -- control passed to block
            Xentry_1386_symbol  <= word_access_1385_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/$entry
            word_access_0_1388: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0 
              signal word_access_0_1388_start: Boolean;
              signal Xentry_1389_symbol: Boolean;
              signal Xexit_1390_symbol: Boolean;
              signal rr_1391_symbol : Boolean;
              signal ra_1392_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1388_start <= Xentry_1386_symbol; -- control passed to block
              Xentry_1389_symbol  <= word_access_0_1388_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/$entry
              rr_1391_symbol <= Xentry_1389_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/rr
              ptr_deref_343_load_0_req_0 <= rr_1391_symbol; -- link to DP
              ra_1392_symbol <= ptr_deref_343_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/ra
              Xexit_1390_symbol <= ra_1392_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0/$exit
              word_access_0_1388_symbol <= Xexit_1390_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/word_access_0
            Xexit_1387_symbol <= word_access_0_1388_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access/$exit
            word_access_1385_symbol <= Xexit_1387_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/word_access
          Xexit_1384_symbol <= word_access_1385_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request/$exit
          ptr_deref_343_request_1382_symbol <= Xexit_1384_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_request
        ptr_deref_343_complete_1393: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete 
          signal ptr_deref_343_complete_1393_start: Boolean;
          signal Xentry_1394_symbol: Boolean;
          signal Xexit_1395_symbol: Boolean;
          signal word_access_1396_symbol : Boolean;
          signal merge_req_1404_symbol : Boolean;
          signal merge_ack_1405_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_343_complete_1393_start <= ptr_deref_343_active_x_x1378_symbol; -- control passed to block
          Xentry_1394_symbol  <= ptr_deref_343_complete_1393_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/$entry
          word_access_1396: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access 
            signal word_access_1396_start: Boolean;
            signal Xentry_1397_symbol: Boolean;
            signal Xexit_1398_symbol: Boolean;
            signal word_access_0_1399_symbol : Boolean;
            -- 
          begin -- 
            word_access_1396_start <= Xentry_1394_symbol; -- control passed to block
            Xentry_1397_symbol  <= word_access_1396_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/$entry
            word_access_0_1399: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0 
              signal word_access_0_1399_start: Boolean;
              signal Xentry_1400_symbol: Boolean;
              signal Xexit_1401_symbol: Boolean;
              signal cr_1402_symbol : Boolean;
              signal ca_1403_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1399_start <= Xentry_1397_symbol; -- control passed to block
              Xentry_1400_symbol  <= word_access_0_1399_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/$entry
              cr_1402_symbol <= Xentry_1400_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/cr
              ptr_deref_343_load_0_req_1 <= cr_1402_symbol; -- link to DP
              ca_1403_symbol <= ptr_deref_343_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/ca
              Xexit_1401_symbol <= ca_1403_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0/$exit
              word_access_0_1399_symbol <= Xexit_1401_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/word_access_0
            Xexit_1398_symbol <= word_access_0_1399_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access/$exit
            word_access_1396_symbol <= Xexit_1398_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/word_access
          merge_req_1404_symbol <= word_access_1396_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/merge_req
          ptr_deref_343_gather_scatter_req_0 <= merge_req_1404_symbol; -- link to DP
          merge_ack_1405_symbol <= ptr_deref_343_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/merge_ack
          Xexit_1395_symbol <= merge_ack_1405_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete/$exit
          ptr_deref_343_complete_1393_symbol <= Xexit_1395_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/ptr_deref_343_complete
        assign_stmt_348_active_x_x1406_symbol <= type_cast_347_complete_1411_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_348_active_
        assign_stmt_348_completed_x_x1407_symbol <= assign_stmt_348_active_x_x1406_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_348_completed_
        type_cast_347_active_x_x1408_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_active_ 
          signal type_cast_347_active_x_x1408_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_347_active_x_x1408_predecessors(0) <= type_cast_347_trigger_x_x1409_symbol;
          type_cast_347_active_x_x1408_predecessors(1) <= simple_obj_ref_346_complete_1410_symbol;
          type_cast_347_active_x_x1408_join: join -- 
            port map( -- 
              preds => type_cast_347_active_x_x1408_predecessors,
              symbol_out => type_cast_347_active_x_x1408_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_active_
        type_cast_347_trigger_x_x1409_symbol <= Xentry_1373_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_trigger_
        simple_obj_ref_346_complete_1410_symbol <= assign_stmt_344_completed_x_x1376_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/simple_obj_ref_346_complete
        type_cast_347_complete_1411: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete 
          signal type_cast_347_complete_1411_start: Boolean;
          signal Xentry_1412_symbol: Boolean;
          signal Xexit_1413_symbol: Boolean;
          signal req_1414_symbol : Boolean;
          signal ack_1415_symbol : Boolean;
          -- 
        begin -- 
          type_cast_347_complete_1411_start <= type_cast_347_active_x_x1408_symbol; -- control passed to block
          Xentry_1412_symbol  <= type_cast_347_complete_1411_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/$entry
          req_1414_symbol <= Xentry_1412_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/req
          type_cast_347_inst_req_0 <= req_1414_symbol; -- link to DP
          ack_1415_symbol <= type_cast_347_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/ack
          Xexit_1413_symbol <= ack_1415_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete/$exit
          type_cast_347_complete_1411_symbol <= Xexit_1413_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/type_cast_347_complete
        assign_stmt_353_active_x_x1416_symbol <= binary_352_complete_1421_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_353_active_
        assign_stmt_353_completed_x_x1417_symbol <= assign_stmt_353_active_x_x1416_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/assign_stmt_353_completed_
        binary_352_active_x_x1418_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_active_ 
          signal binary_352_active_x_x1418_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_352_active_x_x1418_predecessors(0) <= binary_352_trigger_x_x1419_symbol;
          binary_352_active_x_x1418_predecessors(1) <= simple_obj_ref_350_complete_1420_symbol;
          binary_352_active_x_x1418_join: join -- 
            port map( -- 
              preds => binary_352_active_x_x1418_predecessors,
              symbol_out => binary_352_active_x_x1418_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_active_
        binary_352_trigger_x_x1419_symbol <= Xentry_1373_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_trigger_
        simple_obj_ref_350_complete_1420_symbol <= assign_stmt_348_completed_x_x1407_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/simple_obj_ref_350_complete
        binary_352_complete_1421: Block -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete 
          signal binary_352_complete_1421_start: Boolean;
          signal Xentry_1422_symbol: Boolean;
          signal Xexit_1423_symbol: Boolean;
          signal rr_1424_symbol : Boolean;
          signal ra_1425_symbol : Boolean;
          signal cr_1426_symbol : Boolean;
          signal ca_1427_symbol : Boolean;
          -- 
        begin -- 
          binary_352_complete_1421_start <= binary_352_active_x_x1418_symbol; -- control passed to block
          Xentry_1422_symbol  <= binary_352_complete_1421_start; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/$entry
          rr_1424_symbol <= Xentry_1422_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/rr
          binary_352_inst_req_0 <= rr_1424_symbol; -- link to DP
          ra_1425_symbol <= binary_352_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/ra
          cr_1426_symbol <= ra_1425_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/cr
          binary_352_inst_req_1 <= cr_1426_symbol; -- link to DP
          ca_1427_symbol <= binary_352_inst_ack_1; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/ca
          Xexit_1423_symbol <= ca_1427_symbol; -- transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete/$exit
          binary_352_complete_1421_symbol <= Xexit_1423_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/binary_352_complete
        Xexit_1374_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/$exit 
          signal Xexit_1374_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_1374_predecessors(0) <= ptr_deref_343_base_address_calculated_1379_symbol;
          Xexit_1374_predecessors(1) <= assign_stmt_353_completed_x_x1417_symbol;
          Xexit_1374_join: join -- 
            port map( -- 
              preds => Xexit_1374_predecessors,
              symbol_out => Xexit_1374_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353/$exit
        assign_stmt_344_to_assign_stmt_353_1372_symbol <= Xexit_1374_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_344_to_assign_stmt_353
      if_stmt_354_dead_link_1428: Block -- branch_block_stmt_134/if_stmt_354_dead_link 
        signal if_stmt_354_dead_link_1428_start: Boolean;
        signal Xentry_1429_symbol: Boolean;
        signal Xexit_1430_symbol: Boolean;
        signal dead_transition_1431_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_dead_link_1428_start <= if_stmt_354_x_xentry_x_xx_x436_symbol; -- control passed to block
        Xentry_1429_symbol  <= if_stmt_354_dead_link_1428_start; -- transition branch_block_stmt_134/if_stmt_354_dead_link/$entry
        dead_transition_1431_symbol <= false;
        Xexit_1430_symbol <= dead_transition_1431_symbol; -- transition branch_block_stmt_134/if_stmt_354_dead_link/$exit
        if_stmt_354_dead_link_1428_symbol <= Xexit_1430_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_dead_link
      if_stmt_354_eval_test_1432: Block -- branch_block_stmt_134/if_stmt_354_eval_test 
        signal if_stmt_354_eval_test_1432_start: Boolean;
        signal Xentry_1433_symbol: Boolean;
        signal Xexit_1434_symbol: Boolean;
        signal branch_req_1435_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_eval_test_1432_start <= if_stmt_354_x_xentry_x_xx_x436_symbol; -- control passed to block
        Xentry_1433_symbol  <= if_stmt_354_eval_test_1432_start; -- transition branch_block_stmt_134/if_stmt_354_eval_test/$entry
        branch_req_1435_symbol <= Xentry_1433_symbol; -- transition branch_block_stmt_134/if_stmt_354_eval_test/branch_req
        if_stmt_354_branch_req_0 <= branch_req_1435_symbol; -- link to DP
        Xexit_1434_symbol <= branch_req_1435_symbol; -- transition branch_block_stmt_134/if_stmt_354_eval_test/$exit
        if_stmt_354_eval_test_1432_symbol <= Xexit_1434_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_eval_test
      simple_obj_ref_355_place_1436_symbol  <=  if_stmt_354_eval_test_1432_symbol; -- place branch_block_stmt_134/simple_obj_ref_355_place (optimized away) 
      if_stmt_354_if_link_1437: Block -- branch_block_stmt_134/if_stmt_354_if_link 
        signal if_stmt_354_if_link_1437_start: Boolean;
        signal Xentry_1438_symbol: Boolean;
        signal Xexit_1439_symbol: Boolean;
        signal if_choice_transition_1440_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_if_link_1437_start <= simple_obj_ref_355_place_1436_symbol; -- control passed to block
        Xentry_1438_symbol  <= if_stmt_354_if_link_1437_start; -- transition branch_block_stmt_134/if_stmt_354_if_link/$entry
        if_choice_transition_1440_symbol <= if_stmt_354_branch_ack_1; -- transition branch_block_stmt_134/if_stmt_354_if_link/if_choice_transition
        Xexit_1439_symbol <= if_choice_transition_1440_symbol; -- transition branch_block_stmt_134/if_stmt_354_if_link/$exit
        if_stmt_354_if_link_1437_symbol <= Xexit_1439_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_if_link
      if_stmt_354_else_link_1441: Block -- branch_block_stmt_134/if_stmt_354_else_link 
        signal if_stmt_354_else_link_1441_start: Boolean;
        signal Xentry_1442_symbol: Boolean;
        signal Xexit_1443_symbol: Boolean;
        signal else_choice_transition_1444_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_354_else_link_1441_start <= simple_obj_ref_355_place_1436_symbol; -- control passed to block
        Xentry_1442_symbol  <= if_stmt_354_else_link_1441_start; -- transition branch_block_stmt_134/if_stmt_354_else_link/$entry
        else_choice_transition_1444_symbol <= if_stmt_354_branch_ack_0; -- transition branch_block_stmt_134/if_stmt_354_else_link/else_choice_transition
        Xexit_1443_symbol <= else_choice_transition_1444_symbol; -- transition branch_block_stmt_134/if_stmt_354_else_link/$exit
        if_stmt_354_else_link_1441_symbol <= Xexit_1443_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/if_stmt_354_else_link
      bb_8_bb_9_1445_symbol  <=  if_stmt_354_if_link_1437_symbol; -- place branch_block_stmt_134/bb_8_bb_9 (optimized away) 
      bb_8_bb_4_1446_symbol  <=  if_stmt_354_else_link_1441_symbol; -- place branch_block_stmt_134/bb_8_bb_4 (optimized away) 
      assign_stmt_365_1447: Block -- branch_block_stmt_134/assign_stmt_365 
        signal assign_stmt_365_1447_start: Boolean;
        signal Xentry_1448_symbol: Boolean;
        signal Xexit_1449_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_365_1447_start <= assign_stmt_365_x_xentry_x_xx_x440_symbol; -- control passed to block
        Xentry_1448_symbol  <= assign_stmt_365_1447_start; -- transition branch_block_stmt_134/assign_stmt_365/$entry
        Xexit_1449_symbol <= Xentry_1448_symbol; -- transition branch_block_stmt_134/assign_stmt_365/$exit
        assign_stmt_365_1447_symbol <= Xexit_1449_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_365
      assign_stmt_369_1450: Block -- branch_block_stmt_134/assign_stmt_369 
        signal assign_stmt_369_1450_start: Boolean;
        signal Xentry_1451_symbol: Boolean;
        signal Xexit_1452_symbol: Boolean;
        signal assign_stmt_369_active_x_x1453_symbol : Boolean;
        signal assign_stmt_369_completed_x_x1454_symbol : Boolean;
        signal type_cast_368_active_x_x1455_symbol : Boolean;
        signal type_cast_368_trigger_x_x1456_symbol : Boolean;
        signal simple_obj_ref_367_trigger_x_x1457_symbol : Boolean;
        signal simple_obj_ref_367_complete_1458_symbol : Boolean;
        signal type_cast_368_complete_1463_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_369_1450_start <= assign_stmt_369_x_xentry_x_xx_x442_symbol; -- control passed to block
        Xentry_1451_symbol  <= assign_stmt_369_1450_start; -- transition branch_block_stmt_134/assign_stmt_369/$entry
        assign_stmt_369_active_x_x1453_symbol <= type_cast_368_complete_1463_symbol; -- transition branch_block_stmt_134/assign_stmt_369/assign_stmt_369_active_
        assign_stmt_369_completed_x_x1454_symbol <= assign_stmt_369_active_x_x1453_symbol; -- transition branch_block_stmt_134/assign_stmt_369/assign_stmt_369_completed_
        type_cast_368_active_x_x1455_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_369/type_cast_368_active_ 
          signal type_cast_368_active_x_x1455_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_368_active_x_x1455_predecessors(0) <= type_cast_368_trigger_x_x1456_symbol;
          type_cast_368_active_x_x1455_predecessors(1) <= simple_obj_ref_367_complete_1458_symbol;
          type_cast_368_active_x_x1455_join: join -- 
            port map( -- 
              preds => type_cast_368_active_x_x1455_predecessors,
              symbol_out => type_cast_368_active_x_x1455_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_369/type_cast_368_active_
        type_cast_368_trigger_x_x1456_symbol <= Xentry_1451_symbol; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_trigger_
        simple_obj_ref_367_trigger_x_x1457_symbol <= Xentry_1451_symbol; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_trigger_
        simple_obj_ref_367_complete_1458: Block -- branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete 
          signal simple_obj_ref_367_complete_1458_start: Boolean;
          signal Xentry_1459_symbol: Boolean;
          signal Xexit_1460_symbol: Boolean;
          signal req_1461_symbol : Boolean;
          signal ack_1462_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_367_complete_1458_start <= simple_obj_ref_367_trigger_x_x1457_symbol; -- control passed to block
          Xentry_1459_symbol  <= simple_obj_ref_367_complete_1458_start; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/$entry
          req_1461_symbol <= Xentry_1459_symbol; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/req
          simple_obj_ref_367_inst_req_0 <= req_1461_symbol; -- link to DP
          ack_1462_symbol <= simple_obj_ref_367_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/ack
          Xexit_1460_symbol <= ack_1462_symbol; -- transition branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete/$exit
          simple_obj_ref_367_complete_1458_symbol <= Xexit_1460_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_369/simple_obj_ref_367_complete
        type_cast_368_complete_1463: Block -- branch_block_stmt_134/assign_stmt_369/type_cast_368_complete 
          signal type_cast_368_complete_1463_start: Boolean;
          signal Xentry_1464_symbol: Boolean;
          signal Xexit_1465_symbol: Boolean;
          signal req_1466_symbol : Boolean;
          signal ack_1467_symbol : Boolean;
          -- 
        begin -- 
          type_cast_368_complete_1463_start <= type_cast_368_active_x_x1455_symbol; -- control passed to block
          Xentry_1464_symbol  <= type_cast_368_complete_1463_start; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/$entry
          req_1466_symbol <= Xentry_1464_symbol; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/req
          type_cast_368_inst_req_0 <= req_1466_symbol; -- link to DP
          ack_1467_symbol <= type_cast_368_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/ack
          Xexit_1465_symbol <= ack_1467_symbol; -- transition branch_block_stmt_134/assign_stmt_369/type_cast_368_complete/$exit
          type_cast_368_complete_1463_symbol <= Xexit_1465_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_369/type_cast_368_complete
        Xexit_1452_symbol <= assign_stmt_369_completed_x_x1454_symbol; -- transition branch_block_stmt_134/assign_stmt_369/$exit
        assign_stmt_369_1450_symbol <= Xexit_1452_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_369
      assign_stmt_373_to_assign_stmt_400_1468: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400 
        signal assign_stmt_373_to_assign_stmt_400_1468_start: Boolean;
        signal Xentry_1469_symbol: Boolean;
        signal Xexit_1470_symbol: Boolean;
        signal assign_stmt_373_active_x_x1471_symbol : Boolean;
        signal assign_stmt_373_completed_x_x1472_symbol : Boolean;
        signal type_cast_372_active_x_x1473_symbol : Boolean;
        signal type_cast_372_trigger_x_x1474_symbol : Boolean;
        signal simple_obj_ref_371_complete_1475_symbol : Boolean;
        signal type_cast_372_complete_1476_symbol : Boolean;
        signal assign_stmt_377_active_x_x1481_symbol : Boolean;
        signal assign_stmt_377_completed_x_x1482_symbol : Boolean;
        signal simple_obj_ref_376_complete_1483_symbol : Boolean;
        signal ptr_deref_375_trigger_x_x1484_symbol : Boolean;
        signal ptr_deref_375_active_x_x1485_symbol : Boolean;
        signal ptr_deref_375_base_address_calculated_1486_symbol : Boolean;
        signal ptr_deref_375_root_address_calculated_1487_symbol : Boolean;
        signal ptr_deref_375_word_address_calculated_1488_symbol : Boolean;
        signal ptr_deref_375_request_1489_symbol : Boolean;
        signal ptr_deref_375_complete_1502_symbol : Boolean;
        signal assign_stmt_380_active_x_x1513_symbol : Boolean;
        signal assign_stmt_380_completed_x_x1514_symbol : Boolean;
        signal simple_obj_ref_379_trigger_x_x1515_symbol : Boolean;
        signal simple_obj_ref_379_active_x_x1516_symbol : Boolean;
        signal simple_obj_ref_379_root_address_calculated_1517_symbol : Boolean;
        signal simple_obj_ref_379_word_address_calculated_1518_symbol : Boolean;
        signal simple_obj_ref_379_request_1519_symbol : Boolean;
        signal simple_obj_ref_379_complete_1530_symbol : Boolean;
        signal assign_stmt_384_active_x_x1543_symbol : Boolean;
        signal assign_stmt_384_completed_x_x1544_symbol : Boolean;
        signal ptr_deref_383_trigger_x_x1545_symbol : Boolean;
        signal ptr_deref_383_active_x_x1546_symbol : Boolean;
        signal ptr_deref_383_base_address_calculated_1547_symbol : Boolean;
        signal ptr_deref_383_root_address_calculated_1548_symbol : Boolean;
        signal ptr_deref_383_word_address_calculated_1549_symbol : Boolean;
        signal ptr_deref_383_request_1550_symbol : Boolean;
        signal ptr_deref_383_complete_1561_symbol : Boolean;
        signal assign_stmt_389_active_x_x1574_symbol : Boolean;
        signal assign_stmt_389_completed_x_x1575_symbol : Boolean;
        signal array_obj_ref_388_trigger_x_x1576_symbol : Boolean;
        signal array_obj_ref_388_active_x_x1577_symbol : Boolean;
        signal array_obj_ref_388_base_address_calculated_1578_symbol : Boolean;
        signal array_obj_ref_388_root_address_calculated_1579_symbol : Boolean;
        signal array_obj_ref_388_base_address_resized_1580_symbol : Boolean;
        signal array_obj_ref_388_base_addr_resize_1581_symbol : Boolean;
        signal array_obj_ref_388_base_plus_offset_1586_symbol : Boolean;
        signal array_obj_ref_388_complete_1591_symbol : Boolean;
        signal assign_stmt_393_active_x_x1596_symbol : Boolean;
        signal assign_stmt_393_completed_x_x1597_symbol : Boolean;
        signal simple_obj_ref_392_complete_1598_symbol : Boolean;
        signal ptr_deref_391_trigger_x_x1599_symbol : Boolean;
        signal ptr_deref_391_active_x_x1600_symbol : Boolean;
        signal ptr_deref_391_base_address_calculated_1601_symbol : Boolean;
        signal simple_obj_ref_390_complete_1602_symbol : Boolean;
        signal ptr_deref_391_root_address_calculated_1603_symbol : Boolean;
        signal ptr_deref_391_word_address_calculated_1604_symbol : Boolean;
        signal ptr_deref_391_base_address_resized_1605_symbol : Boolean;
        signal ptr_deref_391_base_addr_resize_1606_symbol : Boolean;
        signal ptr_deref_391_base_plus_offset_1611_symbol : Boolean;
        signal ptr_deref_391_word_addrgen_1616_symbol : Boolean;
        signal ptr_deref_391_request_1621_symbol : Boolean;
        signal ptr_deref_391_complete_1634_symbol : Boolean;
        signal assign_stmt_397_active_x_x1645_symbol : Boolean;
        signal assign_stmt_397_completed_x_x1646_symbol : Boolean;
        signal ptr_deref_396_trigger_x_x1647_symbol : Boolean;
        signal ptr_deref_396_active_x_x1648_symbol : Boolean;
        signal ptr_deref_396_base_address_calculated_1649_symbol : Boolean;
        signal ptr_deref_396_root_address_calculated_1650_symbol : Boolean;
        signal ptr_deref_396_word_address_calculated_1651_symbol : Boolean;
        signal ptr_deref_396_request_1652_symbol : Boolean;
        signal ptr_deref_396_complete_1663_symbol : Boolean;
        signal assign_stmt_400_active_x_x1676_symbol : Boolean;
        signal assign_stmt_400_completed_x_x1677_symbol : Boolean;
        signal simple_obj_ref_399_complete_1678_symbol : Boolean;
        signal simple_obj_ref_398_trigger_x_x1679_symbol : Boolean;
        signal simple_obj_ref_398_active_x_x1680_symbol : Boolean;
        signal simple_obj_ref_398_root_address_calculated_1681_symbol : Boolean;
        signal simple_obj_ref_398_word_address_calculated_1682_symbol : Boolean;
        signal simple_obj_ref_398_request_1683_symbol : Boolean;
        signal simple_obj_ref_398_complete_1696_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_373_to_assign_stmt_400_1468_start <= assign_stmt_373_to_assign_stmt_400_x_xentry_x_xx_x444_symbol; -- control passed to block
        Xentry_1469_symbol  <= assign_stmt_373_to_assign_stmt_400_1468_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/$entry
        assign_stmt_373_active_x_x1471_symbol <= type_cast_372_complete_1476_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_373_active_
        assign_stmt_373_completed_x_x1472_symbol <= assign_stmt_373_active_x_x1471_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_373_completed_
        type_cast_372_active_x_x1473_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_active_ 
          signal type_cast_372_active_x_x1473_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_372_active_x_x1473_predecessors(0) <= type_cast_372_trigger_x_x1474_symbol;
          type_cast_372_active_x_x1473_predecessors(1) <= simple_obj_ref_371_complete_1475_symbol;
          type_cast_372_active_x_x1473_join: join -- 
            port map( -- 
              preds => type_cast_372_active_x_x1473_predecessors,
              symbol_out => type_cast_372_active_x_x1473_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_active_
        type_cast_372_trigger_x_x1474_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_trigger_
        simple_obj_ref_371_complete_1475_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_371_complete
        type_cast_372_complete_1476: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete 
          signal type_cast_372_complete_1476_start: Boolean;
          signal Xentry_1477_symbol: Boolean;
          signal Xexit_1478_symbol: Boolean;
          signal req_1479_symbol : Boolean;
          signal ack_1480_symbol : Boolean;
          -- 
        begin -- 
          type_cast_372_complete_1476_start <= type_cast_372_active_x_x1473_symbol; -- control passed to block
          Xentry_1477_symbol  <= type_cast_372_complete_1476_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/$entry
          req_1479_symbol <= Xentry_1477_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/req
          type_cast_372_inst_req_0 <= req_1479_symbol; -- link to DP
          ack_1480_symbol <= type_cast_372_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/ack
          Xexit_1478_symbol <= ack_1480_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete/$exit
          type_cast_372_complete_1476_symbol <= Xexit_1478_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/type_cast_372_complete
        assign_stmt_377_active_x_x1481_symbol <= simple_obj_ref_376_complete_1483_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_377_active_
        assign_stmt_377_completed_x_x1482_symbol <= ptr_deref_375_complete_1502_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_377_completed_
        simple_obj_ref_376_complete_1483_symbol <= assign_stmt_373_completed_x_x1472_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_376_complete
        ptr_deref_375_trigger_x_x1484_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_trigger_ 
          signal ptr_deref_375_trigger_x_x1484_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_375_trigger_x_x1484_predecessors(0) <= ptr_deref_375_word_address_calculated_1488_symbol;
          ptr_deref_375_trigger_x_x1484_predecessors(1) <= assign_stmt_377_active_x_x1481_symbol;
          ptr_deref_375_trigger_x_x1484_join: join -- 
            port map( -- 
              preds => ptr_deref_375_trigger_x_x1484_predecessors,
              symbol_out => ptr_deref_375_trigger_x_x1484_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_trigger_
        ptr_deref_375_active_x_x1485_symbol <= ptr_deref_375_request_1489_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_active_
        ptr_deref_375_base_address_calculated_1486_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_base_address_calculated
        ptr_deref_375_root_address_calculated_1487_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_root_address_calculated
        ptr_deref_375_word_address_calculated_1488_symbol <= ptr_deref_375_root_address_calculated_1487_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_word_address_calculated
        ptr_deref_375_request_1489: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request 
          signal ptr_deref_375_request_1489_start: Boolean;
          signal Xentry_1490_symbol: Boolean;
          signal Xexit_1491_symbol: Boolean;
          signal split_req_1492_symbol : Boolean;
          signal split_ack_1493_symbol : Boolean;
          signal word_access_1494_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_375_request_1489_start <= ptr_deref_375_trigger_x_x1484_symbol; -- control passed to block
          Xentry_1490_symbol  <= ptr_deref_375_request_1489_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/$entry
          split_req_1492_symbol <= Xentry_1490_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/split_req
          ptr_deref_375_gather_scatter_req_0 <= split_req_1492_symbol; -- link to DP
          split_ack_1493_symbol <= ptr_deref_375_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/split_ack
          word_access_1494: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access 
            signal word_access_1494_start: Boolean;
            signal Xentry_1495_symbol: Boolean;
            signal Xexit_1496_symbol: Boolean;
            signal word_access_0_1497_symbol : Boolean;
            -- 
          begin -- 
            word_access_1494_start <= split_ack_1493_symbol; -- control passed to block
            Xentry_1495_symbol  <= word_access_1494_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/$entry
            word_access_0_1497: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0 
              signal word_access_0_1497_start: Boolean;
              signal Xentry_1498_symbol: Boolean;
              signal Xexit_1499_symbol: Boolean;
              signal rr_1500_symbol : Boolean;
              signal ra_1501_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1497_start <= Xentry_1495_symbol; -- control passed to block
              Xentry_1498_symbol  <= word_access_0_1497_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/$entry
              rr_1500_symbol <= Xentry_1498_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/rr
              ptr_deref_375_store_0_req_0 <= rr_1500_symbol; -- link to DP
              ra_1501_symbol <= ptr_deref_375_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/ra
              Xexit_1499_symbol <= ra_1501_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0/$exit
              word_access_0_1497_symbol <= Xexit_1499_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/word_access_0
            Xexit_1496_symbol <= word_access_0_1497_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access/$exit
            word_access_1494_symbol <= Xexit_1496_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/word_access
          Xexit_1491_symbol <= word_access_1494_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request/$exit
          ptr_deref_375_request_1489_symbol <= Xexit_1491_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_request
        ptr_deref_375_complete_1502: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete 
          signal ptr_deref_375_complete_1502_start: Boolean;
          signal Xentry_1503_symbol: Boolean;
          signal Xexit_1504_symbol: Boolean;
          signal word_access_1505_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_375_complete_1502_start <= ptr_deref_375_active_x_x1485_symbol; -- control passed to block
          Xentry_1503_symbol  <= ptr_deref_375_complete_1502_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/$entry
          word_access_1505: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access 
            signal word_access_1505_start: Boolean;
            signal Xentry_1506_symbol: Boolean;
            signal Xexit_1507_symbol: Boolean;
            signal word_access_0_1508_symbol : Boolean;
            -- 
          begin -- 
            word_access_1505_start <= Xentry_1503_symbol; -- control passed to block
            Xentry_1506_symbol  <= word_access_1505_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/$entry
            word_access_0_1508: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0 
              signal word_access_0_1508_start: Boolean;
              signal Xentry_1509_symbol: Boolean;
              signal Xexit_1510_symbol: Boolean;
              signal cr_1511_symbol : Boolean;
              signal ca_1512_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1508_start <= Xentry_1506_symbol; -- control passed to block
              Xentry_1509_symbol  <= word_access_0_1508_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/$entry
              cr_1511_symbol <= Xentry_1509_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/cr
              ptr_deref_375_store_0_req_1 <= cr_1511_symbol; -- link to DP
              ca_1512_symbol <= ptr_deref_375_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/ca
              Xexit_1510_symbol <= ca_1512_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0/$exit
              word_access_0_1508_symbol <= Xexit_1510_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/word_access_0
            Xexit_1507_symbol <= word_access_0_1508_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access/$exit
            word_access_1505_symbol <= Xexit_1507_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/word_access
          Xexit_1504_symbol <= word_access_1505_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete/$exit
          ptr_deref_375_complete_1502_symbol <= Xexit_1504_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_375_complete
        assign_stmt_380_active_x_x1513_symbol <= simple_obj_ref_379_complete_1530_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_380_active_
        assign_stmt_380_completed_x_x1514_symbol <= assign_stmt_380_active_x_x1513_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_380_completed_
        simple_obj_ref_379_trigger_x_x1515_symbol <= simple_obj_ref_379_word_address_calculated_1518_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_trigger_
        simple_obj_ref_379_active_x_x1516_symbol <= simple_obj_ref_379_request_1519_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_active_
        simple_obj_ref_379_root_address_calculated_1517_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_root_address_calculated
        simple_obj_ref_379_word_address_calculated_1518_symbol <= simple_obj_ref_379_root_address_calculated_1517_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_word_address_calculated
        simple_obj_ref_379_request_1519: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request 
          signal simple_obj_ref_379_request_1519_start: Boolean;
          signal Xentry_1520_symbol: Boolean;
          signal Xexit_1521_symbol: Boolean;
          signal word_access_1522_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_379_request_1519_start <= simple_obj_ref_379_trigger_x_x1515_symbol; -- control passed to block
          Xentry_1520_symbol  <= simple_obj_ref_379_request_1519_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/$entry
          word_access_1522: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access 
            signal word_access_1522_start: Boolean;
            signal Xentry_1523_symbol: Boolean;
            signal Xexit_1524_symbol: Boolean;
            signal word_access_0_1525_symbol : Boolean;
            -- 
          begin -- 
            word_access_1522_start <= Xentry_1520_symbol; -- control passed to block
            Xentry_1523_symbol  <= word_access_1522_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/$entry
            word_access_0_1525: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0 
              signal word_access_0_1525_start: Boolean;
              signal Xentry_1526_symbol: Boolean;
              signal Xexit_1527_symbol: Boolean;
              signal rr_1528_symbol : Boolean;
              signal ra_1529_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1525_start <= Xentry_1523_symbol; -- control passed to block
              Xentry_1526_symbol  <= word_access_0_1525_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/$entry
              rr_1528_symbol <= Xentry_1526_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/rr
              simple_obj_ref_379_load_0_req_0 <= rr_1528_symbol; -- link to DP
              ra_1529_symbol <= simple_obj_ref_379_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/ra
              Xexit_1527_symbol <= ra_1529_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0/$exit
              word_access_0_1525_symbol <= Xexit_1527_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/word_access_0
            Xexit_1524_symbol <= word_access_0_1525_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access/$exit
            word_access_1522_symbol <= Xexit_1524_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/word_access
          Xexit_1521_symbol <= word_access_1522_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request/$exit
          simple_obj_ref_379_request_1519_symbol <= Xexit_1521_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_request
        simple_obj_ref_379_complete_1530: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete 
          signal simple_obj_ref_379_complete_1530_start: Boolean;
          signal Xentry_1531_symbol: Boolean;
          signal Xexit_1532_symbol: Boolean;
          signal word_access_1533_symbol : Boolean;
          signal merge_req_1541_symbol : Boolean;
          signal merge_ack_1542_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_379_complete_1530_start <= simple_obj_ref_379_active_x_x1516_symbol; -- control passed to block
          Xentry_1531_symbol  <= simple_obj_ref_379_complete_1530_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/$entry
          word_access_1533: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access 
            signal word_access_1533_start: Boolean;
            signal Xentry_1534_symbol: Boolean;
            signal Xexit_1535_symbol: Boolean;
            signal word_access_0_1536_symbol : Boolean;
            -- 
          begin -- 
            word_access_1533_start <= Xentry_1531_symbol; -- control passed to block
            Xentry_1534_symbol  <= word_access_1533_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/$entry
            word_access_0_1536: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0 
              signal word_access_0_1536_start: Boolean;
              signal Xentry_1537_symbol: Boolean;
              signal Xexit_1538_symbol: Boolean;
              signal cr_1539_symbol : Boolean;
              signal ca_1540_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1536_start <= Xentry_1534_symbol; -- control passed to block
              Xentry_1537_symbol  <= word_access_0_1536_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/$entry
              cr_1539_symbol <= Xentry_1537_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/cr
              simple_obj_ref_379_load_0_req_1 <= cr_1539_symbol; -- link to DP
              ca_1540_symbol <= simple_obj_ref_379_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/ca
              Xexit_1538_symbol <= ca_1540_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0/$exit
              word_access_0_1536_symbol <= Xexit_1538_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/word_access_0
            Xexit_1535_symbol <= word_access_0_1536_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access/$exit
            word_access_1533_symbol <= Xexit_1535_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/word_access
          merge_req_1541_symbol <= word_access_1533_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/merge_req
          simple_obj_ref_379_gather_scatter_req_0 <= merge_req_1541_symbol; -- link to DP
          merge_ack_1542_symbol <= simple_obj_ref_379_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/merge_ack
          Xexit_1532_symbol <= merge_ack_1542_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete/$exit
          simple_obj_ref_379_complete_1530_symbol <= Xexit_1532_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_379_complete
        assign_stmt_384_active_x_x1543_symbol <= ptr_deref_383_complete_1561_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_384_active_
        assign_stmt_384_completed_x_x1544_symbol <= assign_stmt_384_active_x_x1543_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_384_completed_
        ptr_deref_383_trigger_x_x1545_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_trigger_ 
          signal ptr_deref_383_trigger_x_x1545_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_383_trigger_x_x1545_predecessors(0) <= ptr_deref_383_word_address_calculated_1549_symbol;
          ptr_deref_383_trigger_x_x1545_predecessors(1) <= ptr_deref_375_active_x_x1485_symbol;
          ptr_deref_383_trigger_x_x1545_join: join -- 
            port map( -- 
              preds => ptr_deref_383_trigger_x_x1545_predecessors,
              symbol_out => ptr_deref_383_trigger_x_x1545_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_trigger_
        ptr_deref_383_active_x_x1546_symbol <= ptr_deref_383_request_1550_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_active_
        ptr_deref_383_base_address_calculated_1547_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_base_address_calculated
        ptr_deref_383_root_address_calculated_1548_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_root_address_calculated
        ptr_deref_383_word_address_calculated_1549_symbol <= ptr_deref_383_root_address_calculated_1548_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_word_address_calculated
        ptr_deref_383_request_1550: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request 
          signal ptr_deref_383_request_1550_start: Boolean;
          signal Xentry_1551_symbol: Boolean;
          signal Xexit_1552_symbol: Boolean;
          signal word_access_1553_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_383_request_1550_start <= ptr_deref_383_trigger_x_x1545_symbol; -- control passed to block
          Xentry_1551_symbol  <= ptr_deref_383_request_1550_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/$entry
          word_access_1553: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access 
            signal word_access_1553_start: Boolean;
            signal Xentry_1554_symbol: Boolean;
            signal Xexit_1555_symbol: Boolean;
            signal word_access_0_1556_symbol : Boolean;
            -- 
          begin -- 
            word_access_1553_start <= Xentry_1551_symbol; -- control passed to block
            Xentry_1554_symbol  <= word_access_1553_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/$entry
            word_access_0_1556: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0 
              signal word_access_0_1556_start: Boolean;
              signal Xentry_1557_symbol: Boolean;
              signal Xexit_1558_symbol: Boolean;
              signal rr_1559_symbol : Boolean;
              signal ra_1560_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1556_start <= Xentry_1554_symbol; -- control passed to block
              Xentry_1557_symbol  <= word_access_0_1556_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/$entry
              rr_1559_symbol <= Xentry_1557_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/rr
              ptr_deref_383_load_0_req_0 <= rr_1559_symbol; -- link to DP
              ra_1560_symbol <= ptr_deref_383_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/ra
              Xexit_1558_symbol <= ra_1560_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0/$exit
              word_access_0_1556_symbol <= Xexit_1558_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/word_access_0
            Xexit_1555_symbol <= word_access_0_1556_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access/$exit
            word_access_1553_symbol <= Xexit_1555_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/word_access
          Xexit_1552_symbol <= word_access_1553_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request/$exit
          ptr_deref_383_request_1550_symbol <= Xexit_1552_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_request
        ptr_deref_383_complete_1561: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete 
          signal ptr_deref_383_complete_1561_start: Boolean;
          signal Xentry_1562_symbol: Boolean;
          signal Xexit_1563_symbol: Boolean;
          signal word_access_1564_symbol : Boolean;
          signal merge_req_1572_symbol : Boolean;
          signal merge_ack_1573_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_383_complete_1561_start <= ptr_deref_383_active_x_x1546_symbol; -- control passed to block
          Xentry_1562_symbol  <= ptr_deref_383_complete_1561_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/$entry
          word_access_1564: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access 
            signal word_access_1564_start: Boolean;
            signal Xentry_1565_symbol: Boolean;
            signal Xexit_1566_symbol: Boolean;
            signal word_access_0_1567_symbol : Boolean;
            -- 
          begin -- 
            word_access_1564_start <= Xentry_1562_symbol; -- control passed to block
            Xentry_1565_symbol  <= word_access_1564_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/$entry
            word_access_0_1567: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0 
              signal word_access_0_1567_start: Boolean;
              signal Xentry_1568_symbol: Boolean;
              signal Xexit_1569_symbol: Boolean;
              signal cr_1570_symbol : Boolean;
              signal ca_1571_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1567_start <= Xentry_1565_symbol; -- control passed to block
              Xentry_1568_symbol  <= word_access_0_1567_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/$entry
              cr_1570_symbol <= Xentry_1568_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/cr
              ptr_deref_383_load_0_req_1 <= cr_1570_symbol; -- link to DP
              ca_1571_symbol <= ptr_deref_383_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/ca
              Xexit_1569_symbol <= ca_1571_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0/$exit
              word_access_0_1567_symbol <= Xexit_1569_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/word_access_0
            Xexit_1566_symbol <= word_access_0_1567_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access/$exit
            word_access_1564_symbol <= Xexit_1566_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/word_access
          merge_req_1572_symbol <= word_access_1564_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/merge_req
          ptr_deref_383_gather_scatter_req_0 <= merge_req_1572_symbol; -- link to DP
          merge_ack_1573_symbol <= ptr_deref_383_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/merge_ack
          Xexit_1563_symbol <= merge_ack_1573_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete/$exit
          ptr_deref_383_complete_1561_symbol <= Xexit_1563_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_383_complete
        assign_stmt_389_active_x_x1574_symbol <= array_obj_ref_388_complete_1591_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_389_active_
        assign_stmt_389_completed_x_x1575_symbol <= assign_stmt_389_active_x_x1574_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_389_completed_
        array_obj_ref_388_trigger_x_x1576_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_trigger_
        array_obj_ref_388_active_x_x1577_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_active_ 
          signal array_obj_ref_388_active_x_x1577_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_388_active_x_x1577_predecessors(0) <= array_obj_ref_388_trigger_x_x1576_symbol;
          array_obj_ref_388_active_x_x1577_predecessors(1) <= array_obj_ref_388_root_address_calculated_1579_symbol;
          array_obj_ref_388_active_x_x1577_join: join -- 
            port map( -- 
              preds => array_obj_ref_388_active_x_x1577_predecessors,
              symbol_out => array_obj_ref_388_active_x_x1577_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_active_
        array_obj_ref_388_base_address_calculated_1578_symbol <= assign_stmt_384_completed_x_x1544_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_address_calculated
        array_obj_ref_388_root_address_calculated_1579_symbol <= array_obj_ref_388_base_plus_offset_1586_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_root_address_calculated
        array_obj_ref_388_base_address_resized_1580_symbol <= array_obj_ref_388_base_addr_resize_1581_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_address_resized
        array_obj_ref_388_base_addr_resize_1581: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize 
          signal array_obj_ref_388_base_addr_resize_1581_start: Boolean;
          signal Xentry_1582_symbol: Boolean;
          signal Xexit_1583_symbol: Boolean;
          signal base_resize_req_1584_symbol : Boolean;
          signal base_resize_ack_1585_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_388_base_addr_resize_1581_start <= array_obj_ref_388_base_address_calculated_1578_symbol; -- control passed to block
          Xentry_1582_symbol  <= array_obj_ref_388_base_addr_resize_1581_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/$entry
          base_resize_req_1584_symbol <= Xentry_1582_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/base_resize_req
          array_obj_ref_388_base_resize_req_0 <= base_resize_req_1584_symbol; -- link to DP
          base_resize_ack_1585_symbol <= array_obj_ref_388_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/base_resize_ack
          Xexit_1583_symbol <= base_resize_ack_1585_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize/$exit
          array_obj_ref_388_base_addr_resize_1581_symbol <= Xexit_1583_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_addr_resize
        array_obj_ref_388_base_plus_offset_1586: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset 
          signal array_obj_ref_388_base_plus_offset_1586_start: Boolean;
          signal Xentry_1587_symbol: Boolean;
          signal Xexit_1588_symbol: Boolean;
          signal sum_rename_req_1589_symbol : Boolean;
          signal sum_rename_ack_1590_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_388_base_plus_offset_1586_start <= array_obj_ref_388_base_address_resized_1580_symbol; -- control passed to block
          Xentry_1587_symbol  <= array_obj_ref_388_base_plus_offset_1586_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/$entry
          sum_rename_req_1589_symbol <= Xentry_1587_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/sum_rename_req
          array_obj_ref_388_root_address_inst_req_0 <= sum_rename_req_1589_symbol; -- link to DP
          sum_rename_ack_1590_symbol <= array_obj_ref_388_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/sum_rename_ack
          Xexit_1588_symbol <= sum_rename_ack_1590_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset/$exit
          array_obj_ref_388_base_plus_offset_1586_symbol <= Xexit_1588_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_base_plus_offset
        array_obj_ref_388_complete_1591: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete 
          signal array_obj_ref_388_complete_1591_start: Boolean;
          signal Xentry_1592_symbol: Boolean;
          signal Xexit_1593_symbol: Boolean;
          signal final_reg_req_1594_symbol : Boolean;
          signal final_reg_ack_1595_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_388_complete_1591_start <= array_obj_ref_388_active_x_x1577_symbol; -- control passed to block
          Xentry_1592_symbol  <= array_obj_ref_388_complete_1591_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/$entry
          final_reg_req_1594_symbol <= Xentry_1592_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/final_reg_req
          array_obj_ref_388_final_reg_req_0 <= final_reg_req_1594_symbol; -- link to DP
          final_reg_ack_1595_symbol <= array_obj_ref_388_final_reg_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/final_reg_ack
          Xexit_1593_symbol <= final_reg_ack_1595_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete/$exit
          array_obj_ref_388_complete_1591_symbol <= Xexit_1593_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/array_obj_ref_388_complete
        assign_stmt_393_active_x_x1596_symbol <= simple_obj_ref_392_complete_1598_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_393_active_
        assign_stmt_393_completed_x_x1597_symbol <= ptr_deref_391_complete_1634_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_393_completed_
        simple_obj_ref_392_complete_1598_symbol <= assign_stmt_380_completed_x_x1514_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_392_complete
        ptr_deref_391_trigger_x_x1599_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_trigger_ 
          signal ptr_deref_391_trigger_x_x1599_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          ptr_deref_391_trigger_x_x1599_predecessors(0) <= ptr_deref_391_word_address_calculated_1604_symbol;
          ptr_deref_391_trigger_x_x1599_predecessors(1) <= ptr_deref_391_base_address_calculated_1601_symbol;
          ptr_deref_391_trigger_x_x1599_predecessors(2) <= assign_stmt_393_active_x_x1596_symbol;
          ptr_deref_391_trigger_x_x1599_join: join -- 
            port map( -- 
              preds => ptr_deref_391_trigger_x_x1599_predecessors,
              symbol_out => ptr_deref_391_trigger_x_x1599_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_trigger_
        ptr_deref_391_active_x_x1600_symbol <= ptr_deref_391_request_1621_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_active_
        ptr_deref_391_base_address_calculated_1601_symbol <= simple_obj_ref_390_complete_1602_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_address_calculated
        simple_obj_ref_390_complete_1602_symbol <= assign_stmt_389_completed_x_x1575_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_390_complete
        ptr_deref_391_root_address_calculated_1603_symbol <= ptr_deref_391_base_plus_offset_1611_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_root_address_calculated
        ptr_deref_391_word_address_calculated_1604_symbol <= ptr_deref_391_word_addrgen_1616_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_address_calculated
        ptr_deref_391_base_address_resized_1605_symbol <= ptr_deref_391_base_addr_resize_1606_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_address_resized
        ptr_deref_391_base_addr_resize_1606: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize 
          signal ptr_deref_391_base_addr_resize_1606_start: Boolean;
          signal Xentry_1607_symbol: Boolean;
          signal Xexit_1608_symbol: Boolean;
          signal base_resize_req_1609_symbol : Boolean;
          signal base_resize_ack_1610_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_base_addr_resize_1606_start <= ptr_deref_391_base_address_calculated_1601_symbol; -- control passed to block
          Xentry_1607_symbol  <= ptr_deref_391_base_addr_resize_1606_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/$entry
          base_resize_req_1609_symbol <= Xentry_1607_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/base_resize_req
          ptr_deref_391_base_resize_req_0 <= base_resize_req_1609_symbol; -- link to DP
          base_resize_ack_1610_symbol <= ptr_deref_391_base_resize_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/base_resize_ack
          Xexit_1608_symbol <= base_resize_ack_1610_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize/$exit
          ptr_deref_391_base_addr_resize_1606_symbol <= Xexit_1608_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_addr_resize
        ptr_deref_391_base_plus_offset_1611: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset 
          signal ptr_deref_391_base_plus_offset_1611_start: Boolean;
          signal Xentry_1612_symbol: Boolean;
          signal Xexit_1613_symbol: Boolean;
          signal sum_rename_req_1614_symbol : Boolean;
          signal sum_rename_ack_1615_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_base_plus_offset_1611_start <= ptr_deref_391_base_address_resized_1605_symbol; -- control passed to block
          Xentry_1612_symbol  <= ptr_deref_391_base_plus_offset_1611_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/$entry
          sum_rename_req_1614_symbol <= Xentry_1612_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/sum_rename_req
          ptr_deref_391_root_address_inst_req_0 <= sum_rename_req_1614_symbol; -- link to DP
          sum_rename_ack_1615_symbol <= ptr_deref_391_root_address_inst_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/sum_rename_ack
          Xexit_1613_symbol <= sum_rename_ack_1615_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset/$exit
          ptr_deref_391_base_plus_offset_1611_symbol <= Xexit_1613_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_base_plus_offset
        ptr_deref_391_word_addrgen_1616: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen 
          signal ptr_deref_391_word_addrgen_1616_start: Boolean;
          signal Xentry_1617_symbol: Boolean;
          signal Xexit_1618_symbol: Boolean;
          signal root_rename_req_1619_symbol : Boolean;
          signal root_rename_ack_1620_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_word_addrgen_1616_start <= ptr_deref_391_root_address_calculated_1603_symbol; -- control passed to block
          Xentry_1617_symbol  <= ptr_deref_391_word_addrgen_1616_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/$entry
          root_rename_req_1619_symbol <= Xentry_1617_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/root_rename_req
          ptr_deref_391_addr_0_req_0 <= root_rename_req_1619_symbol; -- link to DP
          root_rename_ack_1620_symbol <= ptr_deref_391_addr_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/root_rename_ack
          Xexit_1618_symbol <= root_rename_ack_1620_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen/$exit
          ptr_deref_391_word_addrgen_1616_symbol <= Xexit_1618_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_word_addrgen
        ptr_deref_391_request_1621: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request 
          signal ptr_deref_391_request_1621_start: Boolean;
          signal Xentry_1622_symbol: Boolean;
          signal Xexit_1623_symbol: Boolean;
          signal split_req_1624_symbol : Boolean;
          signal split_ack_1625_symbol : Boolean;
          signal word_access_1626_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_request_1621_start <= ptr_deref_391_trigger_x_x1599_symbol; -- control passed to block
          Xentry_1622_symbol  <= ptr_deref_391_request_1621_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/$entry
          split_req_1624_symbol <= Xentry_1622_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/split_req
          ptr_deref_391_gather_scatter_req_0 <= split_req_1624_symbol; -- link to DP
          split_ack_1625_symbol <= ptr_deref_391_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/split_ack
          word_access_1626: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access 
            signal word_access_1626_start: Boolean;
            signal Xentry_1627_symbol: Boolean;
            signal Xexit_1628_symbol: Boolean;
            signal word_access_0_1629_symbol : Boolean;
            -- 
          begin -- 
            word_access_1626_start <= split_ack_1625_symbol; -- control passed to block
            Xentry_1627_symbol  <= word_access_1626_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/$entry
            word_access_0_1629: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0 
              signal word_access_0_1629_start: Boolean;
              signal Xentry_1630_symbol: Boolean;
              signal Xexit_1631_symbol: Boolean;
              signal rr_1632_symbol : Boolean;
              signal ra_1633_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1629_start <= Xentry_1627_symbol; -- control passed to block
              Xentry_1630_symbol  <= word_access_0_1629_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/$entry
              rr_1632_symbol <= Xentry_1630_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/rr
              ptr_deref_391_store_0_req_0 <= rr_1632_symbol; -- link to DP
              ra_1633_symbol <= ptr_deref_391_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/ra
              Xexit_1631_symbol <= ra_1633_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0/$exit
              word_access_0_1629_symbol <= Xexit_1631_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/word_access_0
            Xexit_1628_symbol <= word_access_0_1629_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access/$exit
            word_access_1626_symbol <= Xexit_1628_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/word_access
          Xexit_1623_symbol <= word_access_1626_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request/$exit
          ptr_deref_391_request_1621_symbol <= Xexit_1623_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_request
        ptr_deref_391_complete_1634: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete 
          signal ptr_deref_391_complete_1634_start: Boolean;
          signal Xentry_1635_symbol: Boolean;
          signal Xexit_1636_symbol: Boolean;
          signal word_access_1637_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_391_complete_1634_start <= ptr_deref_391_active_x_x1600_symbol; -- control passed to block
          Xentry_1635_symbol  <= ptr_deref_391_complete_1634_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/$entry
          word_access_1637: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access 
            signal word_access_1637_start: Boolean;
            signal Xentry_1638_symbol: Boolean;
            signal Xexit_1639_symbol: Boolean;
            signal word_access_0_1640_symbol : Boolean;
            -- 
          begin -- 
            word_access_1637_start <= Xentry_1635_symbol; -- control passed to block
            Xentry_1638_symbol  <= word_access_1637_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/$entry
            word_access_0_1640: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0 
              signal word_access_0_1640_start: Boolean;
              signal Xentry_1641_symbol: Boolean;
              signal Xexit_1642_symbol: Boolean;
              signal cr_1643_symbol : Boolean;
              signal ca_1644_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1640_start <= Xentry_1638_symbol; -- control passed to block
              Xentry_1641_symbol  <= word_access_0_1640_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/$entry
              cr_1643_symbol <= Xentry_1641_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/cr
              ptr_deref_391_store_0_req_1 <= cr_1643_symbol; -- link to DP
              ca_1644_symbol <= ptr_deref_391_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/ca
              Xexit_1642_symbol <= ca_1644_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0/$exit
              word_access_0_1640_symbol <= Xexit_1642_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/word_access_0
            Xexit_1639_symbol <= word_access_0_1640_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access/$exit
            word_access_1637_symbol <= Xexit_1639_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/word_access
          Xexit_1636_symbol <= word_access_1637_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete/$exit
          ptr_deref_391_complete_1634_symbol <= Xexit_1636_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_391_complete
        assign_stmt_397_active_x_x1645_symbol <= ptr_deref_396_complete_1663_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_397_active_
        assign_stmt_397_completed_x_x1646_symbol <= assign_stmt_397_active_x_x1645_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_397_completed_
        ptr_deref_396_trigger_x_x1647_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_trigger_ 
          signal ptr_deref_396_trigger_x_x1647_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_396_trigger_x_x1647_predecessors(0) <= ptr_deref_396_word_address_calculated_1651_symbol;
          ptr_deref_396_trigger_x_x1647_predecessors(1) <= ptr_deref_375_active_x_x1485_symbol;
          ptr_deref_396_trigger_x_x1647_join: join -- 
            port map( -- 
              preds => ptr_deref_396_trigger_x_x1647_predecessors,
              symbol_out => ptr_deref_396_trigger_x_x1647_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_trigger_
        ptr_deref_396_active_x_x1648_symbol <= ptr_deref_396_request_1652_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_active_
        ptr_deref_396_base_address_calculated_1649_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_base_address_calculated
        ptr_deref_396_root_address_calculated_1650_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_root_address_calculated
        ptr_deref_396_word_address_calculated_1651_symbol <= ptr_deref_396_root_address_calculated_1650_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_word_address_calculated
        ptr_deref_396_request_1652: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request 
          signal ptr_deref_396_request_1652_start: Boolean;
          signal Xentry_1653_symbol: Boolean;
          signal Xexit_1654_symbol: Boolean;
          signal word_access_1655_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_396_request_1652_start <= ptr_deref_396_trigger_x_x1647_symbol; -- control passed to block
          Xentry_1653_symbol  <= ptr_deref_396_request_1652_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/$entry
          word_access_1655: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access 
            signal word_access_1655_start: Boolean;
            signal Xentry_1656_symbol: Boolean;
            signal Xexit_1657_symbol: Boolean;
            signal word_access_0_1658_symbol : Boolean;
            -- 
          begin -- 
            word_access_1655_start <= Xentry_1653_symbol; -- control passed to block
            Xentry_1656_symbol  <= word_access_1655_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/$entry
            word_access_0_1658: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0 
              signal word_access_0_1658_start: Boolean;
              signal Xentry_1659_symbol: Boolean;
              signal Xexit_1660_symbol: Boolean;
              signal rr_1661_symbol : Boolean;
              signal ra_1662_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1658_start <= Xentry_1656_symbol; -- control passed to block
              Xentry_1659_symbol  <= word_access_0_1658_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/$entry
              rr_1661_symbol <= Xentry_1659_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/rr
              ptr_deref_396_load_0_req_0 <= rr_1661_symbol; -- link to DP
              ra_1662_symbol <= ptr_deref_396_load_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/ra
              Xexit_1660_symbol <= ra_1662_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0/$exit
              word_access_0_1658_symbol <= Xexit_1660_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/word_access_0
            Xexit_1657_symbol <= word_access_0_1658_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access/$exit
            word_access_1655_symbol <= Xexit_1657_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/word_access
          Xexit_1654_symbol <= word_access_1655_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request/$exit
          ptr_deref_396_request_1652_symbol <= Xexit_1654_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_request
        ptr_deref_396_complete_1663: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete 
          signal ptr_deref_396_complete_1663_start: Boolean;
          signal Xentry_1664_symbol: Boolean;
          signal Xexit_1665_symbol: Boolean;
          signal word_access_1666_symbol : Boolean;
          signal merge_req_1674_symbol : Boolean;
          signal merge_ack_1675_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_396_complete_1663_start <= ptr_deref_396_active_x_x1648_symbol; -- control passed to block
          Xentry_1664_symbol  <= ptr_deref_396_complete_1663_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/$entry
          word_access_1666: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access 
            signal word_access_1666_start: Boolean;
            signal Xentry_1667_symbol: Boolean;
            signal Xexit_1668_symbol: Boolean;
            signal word_access_0_1669_symbol : Boolean;
            -- 
          begin -- 
            word_access_1666_start <= Xentry_1664_symbol; -- control passed to block
            Xentry_1667_symbol  <= word_access_1666_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/$entry
            word_access_0_1669: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0 
              signal word_access_0_1669_start: Boolean;
              signal Xentry_1670_symbol: Boolean;
              signal Xexit_1671_symbol: Boolean;
              signal cr_1672_symbol : Boolean;
              signal ca_1673_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1669_start <= Xentry_1667_symbol; -- control passed to block
              Xentry_1670_symbol  <= word_access_0_1669_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/$entry
              cr_1672_symbol <= Xentry_1670_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/cr
              ptr_deref_396_load_0_req_1 <= cr_1672_symbol; -- link to DP
              ca_1673_symbol <= ptr_deref_396_load_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/ca
              Xexit_1671_symbol <= ca_1673_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0/$exit
              word_access_0_1669_symbol <= Xexit_1671_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/word_access_0
            Xexit_1668_symbol <= word_access_0_1669_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access/$exit
            word_access_1666_symbol <= Xexit_1668_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/word_access
          merge_req_1674_symbol <= word_access_1666_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/merge_req
          ptr_deref_396_gather_scatter_req_0 <= merge_req_1674_symbol; -- link to DP
          merge_ack_1675_symbol <= ptr_deref_396_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/merge_ack
          Xexit_1665_symbol <= merge_ack_1675_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete/$exit
          ptr_deref_396_complete_1663_symbol <= Xexit_1665_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/ptr_deref_396_complete
        assign_stmt_400_active_x_x1676_symbol <= simple_obj_ref_399_complete_1678_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_400_active_
        assign_stmt_400_completed_x_x1677_symbol <= simple_obj_ref_398_complete_1696_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/assign_stmt_400_completed_
        simple_obj_ref_399_complete_1678_symbol <= assign_stmt_397_completed_x_x1646_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_399_complete
        simple_obj_ref_398_trigger_x_x1679_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_trigger_ 
          signal simple_obj_ref_398_trigger_x_x1679_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          simple_obj_ref_398_trigger_x_x1679_predecessors(0) <= simple_obj_ref_398_word_address_calculated_1682_symbol;
          simple_obj_ref_398_trigger_x_x1679_predecessors(1) <= assign_stmt_400_active_x_x1676_symbol;
          simple_obj_ref_398_trigger_x_x1679_predecessors(2) <= simple_obj_ref_379_active_x_x1516_symbol;
          simple_obj_ref_398_trigger_x_x1679_join: join -- 
            port map( -- 
              preds => simple_obj_ref_398_trigger_x_x1679_predecessors,
              symbol_out => simple_obj_ref_398_trigger_x_x1679_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_trigger_
        simple_obj_ref_398_active_x_x1680_symbol <= simple_obj_ref_398_request_1683_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_active_
        simple_obj_ref_398_root_address_calculated_1681_symbol <= Xentry_1469_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_root_address_calculated
        simple_obj_ref_398_word_address_calculated_1682_symbol <= simple_obj_ref_398_root_address_calculated_1681_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_word_address_calculated
        simple_obj_ref_398_request_1683: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request 
          signal simple_obj_ref_398_request_1683_start: Boolean;
          signal Xentry_1684_symbol: Boolean;
          signal Xexit_1685_symbol: Boolean;
          signal split_req_1686_symbol : Boolean;
          signal split_ack_1687_symbol : Boolean;
          signal word_access_1688_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_398_request_1683_start <= simple_obj_ref_398_trigger_x_x1679_symbol; -- control passed to block
          Xentry_1684_symbol  <= simple_obj_ref_398_request_1683_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/$entry
          split_req_1686_symbol <= Xentry_1684_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/split_req
          simple_obj_ref_398_gather_scatter_req_0 <= split_req_1686_symbol; -- link to DP
          split_ack_1687_symbol <= simple_obj_ref_398_gather_scatter_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/split_ack
          word_access_1688: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access 
            signal word_access_1688_start: Boolean;
            signal Xentry_1689_symbol: Boolean;
            signal Xexit_1690_symbol: Boolean;
            signal word_access_0_1691_symbol : Boolean;
            -- 
          begin -- 
            word_access_1688_start <= split_ack_1687_symbol; -- control passed to block
            Xentry_1689_symbol  <= word_access_1688_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/$entry
            word_access_0_1691: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0 
              signal word_access_0_1691_start: Boolean;
              signal Xentry_1692_symbol: Boolean;
              signal Xexit_1693_symbol: Boolean;
              signal rr_1694_symbol : Boolean;
              signal ra_1695_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1691_start <= Xentry_1689_symbol; -- control passed to block
              Xentry_1692_symbol  <= word_access_0_1691_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/$entry
              rr_1694_symbol <= Xentry_1692_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/rr
              simple_obj_ref_398_store_0_req_0 <= rr_1694_symbol; -- link to DP
              ra_1695_symbol <= simple_obj_ref_398_store_0_ack_0; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/ra
              Xexit_1693_symbol <= ra_1695_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0/$exit
              word_access_0_1691_symbol <= Xexit_1693_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/word_access_0
            Xexit_1690_symbol <= word_access_0_1691_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access/$exit
            word_access_1688_symbol <= Xexit_1690_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/word_access
          Xexit_1685_symbol <= word_access_1688_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request/$exit
          simple_obj_ref_398_request_1683_symbol <= Xexit_1685_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_request
        simple_obj_ref_398_complete_1696: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete 
          signal simple_obj_ref_398_complete_1696_start: Boolean;
          signal Xentry_1697_symbol: Boolean;
          signal Xexit_1698_symbol: Boolean;
          signal word_access_1699_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_398_complete_1696_start <= simple_obj_ref_398_active_x_x1680_symbol; -- control passed to block
          Xentry_1697_symbol  <= simple_obj_ref_398_complete_1696_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/$entry
          word_access_1699: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access 
            signal word_access_1699_start: Boolean;
            signal Xentry_1700_symbol: Boolean;
            signal Xexit_1701_symbol: Boolean;
            signal word_access_0_1702_symbol : Boolean;
            -- 
          begin -- 
            word_access_1699_start <= Xentry_1697_symbol; -- control passed to block
            Xentry_1700_symbol  <= word_access_1699_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/$entry
            word_access_0_1702: Block -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0 
              signal word_access_0_1702_start: Boolean;
              signal Xentry_1703_symbol: Boolean;
              signal Xexit_1704_symbol: Boolean;
              signal cr_1705_symbol : Boolean;
              signal ca_1706_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1702_start <= Xentry_1700_symbol; -- control passed to block
              Xentry_1703_symbol  <= word_access_0_1702_start; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/$entry
              cr_1705_symbol <= Xentry_1703_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/cr
              simple_obj_ref_398_store_0_req_1 <= cr_1705_symbol; -- link to DP
              ca_1706_symbol <= simple_obj_ref_398_store_0_ack_1; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/ca
              Xexit_1704_symbol <= ca_1706_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0/$exit
              word_access_0_1702_symbol <= Xexit_1704_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/word_access_0
            Xexit_1701_symbol <= word_access_0_1702_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access/$exit
            word_access_1699_symbol <= Xexit_1701_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/word_access
          Xexit_1698_symbol <= word_access_1699_symbol; -- transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete/$exit
          simple_obj_ref_398_complete_1696_symbol <= Xexit_1698_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/simple_obj_ref_398_complete
        Xexit_1470_block : Block -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/$exit 
          signal Xexit_1470_predecessors: BooleanArray(5 downto 0);
          -- 
        begin -- 
          Xexit_1470_predecessors(0) <= assign_stmt_377_completed_x_x1482_symbol;
          Xexit_1470_predecessors(1) <= ptr_deref_375_base_address_calculated_1486_symbol;
          Xexit_1470_predecessors(2) <= ptr_deref_383_base_address_calculated_1547_symbol;
          Xexit_1470_predecessors(3) <= assign_stmt_393_completed_x_x1597_symbol;
          Xexit_1470_predecessors(4) <= ptr_deref_396_base_address_calculated_1649_symbol;
          Xexit_1470_predecessors(5) <= assign_stmt_400_completed_x_x1677_symbol;
          Xexit_1470_join: join -- 
            port map( -- 
              preds => Xexit_1470_predecessors,
              symbol_out => Xexit_1470_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400/$exit
        assign_stmt_373_to_assign_stmt_400_1468_symbol <= Xexit_1470_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/assign_stmt_373_to_assign_stmt_400
      bb_0_bb_1_PhiReq_1707: Block -- branch_block_stmt_134/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_1707_start: Boolean;
        signal Xentry_1708_symbol: Boolean;
        signal Xexit_1709_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_1707_start <= bb_0_bb_1_392_symbol; -- control passed to block
        Xentry_1708_symbol  <= bb_0_bb_1_PhiReq_1707_start; -- transition branch_block_stmt_134/bb_0_bb_1_PhiReq/$entry
        Xexit_1709_symbol <= Xentry_1708_symbol; -- transition branch_block_stmt_134/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_1707_symbol <= Xexit_1709_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_0_bb_1_PhiReq
      bb_2_bb_1_PhiReq_1710: Block -- branch_block_stmt_134/bb_2_bb_1_PhiReq 
        signal bb_2_bb_1_PhiReq_1710_start: Boolean;
        signal Xentry_1711_symbol: Boolean;
        signal Xexit_1712_symbol: Boolean;
        -- 
      begin -- 
        bb_2_bb_1_PhiReq_1710_start <= bb_2_bb_1_402_symbol; -- control passed to block
        Xentry_1711_symbol  <= bb_2_bb_1_PhiReq_1710_start; -- transition branch_block_stmt_134/bb_2_bb_1_PhiReq/$entry
        Xexit_1712_symbol <= Xentry_1711_symbol; -- transition branch_block_stmt_134/bb_2_bb_1_PhiReq/$exit
        bb_2_bb_1_PhiReq_1710_symbol <= Xexit_1712_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_2_bb_1_PhiReq
      merge_stmt_160_PhiReqMerge_1713_symbol  <=  bb_0_bb_1_PhiReq_1707_symbol or bb_2_bb_1_PhiReq_1710_symbol; -- place branch_block_stmt_134/merge_stmt_160_PhiReqMerge (optimized away) 
      merge_stmt_160_PhiAck_1714: Block -- branch_block_stmt_134/merge_stmt_160_PhiAck 
        signal merge_stmt_160_PhiAck_1714_start: Boolean;
        signal Xentry_1715_symbol: Boolean;
        signal Xexit_1716_symbol: Boolean;
        signal dummy_1717_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_160_PhiAck_1714_start <= merge_stmt_160_PhiReqMerge_1713_symbol; -- control passed to block
        Xentry_1715_symbol  <= merge_stmt_160_PhiAck_1714_start; -- transition branch_block_stmt_134/merge_stmt_160_PhiAck/$entry
        dummy_1717_symbol <= Xentry_1715_symbol; -- transition branch_block_stmt_134/merge_stmt_160_PhiAck/dummy
        Xexit_1716_symbol <= dummy_1717_symbol; -- transition branch_block_stmt_134/merge_stmt_160_PhiAck/$exit
        merge_stmt_160_PhiAck_1714_symbol <= Xexit_1716_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_160_PhiAck
      merge_stmt_180_dead_link_1718: Block -- branch_block_stmt_134/merge_stmt_180_dead_link 
        signal merge_stmt_180_dead_link_1718_start: Boolean;
        signal Xentry_1719_symbol: Boolean;
        signal Xexit_1720_symbol: Boolean;
        signal dead_transition_1721_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_180_dead_link_1718_start <= merge_stmt_180_x_xentry_x_xx_x398_symbol; -- control passed to block
        Xentry_1719_symbol  <= merge_stmt_180_dead_link_1718_start; -- transition branch_block_stmt_134/merge_stmt_180_dead_link/$entry
        dead_transition_1721_symbol <= false;
        Xexit_1720_symbol <= dead_transition_1721_symbol; -- transition branch_block_stmt_134/merge_stmt_180_dead_link/$exit
        merge_stmt_180_dead_link_1718_symbol <= Xexit_1720_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_180_dead_link
      bb_1_bb_2_PhiReq_1722: Block -- branch_block_stmt_134/bb_1_bb_2_PhiReq 
        signal bb_1_bb_2_PhiReq_1722_start: Boolean;
        signal Xentry_1723_symbol: Boolean;
        signal Xexit_1724_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_2_PhiReq_1722_start <= bb_1_bb_2_551_symbol; -- control passed to block
        Xentry_1723_symbol  <= bb_1_bb_2_PhiReq_1722_start; -- transition branch_block_stmt_134/bb_1_bb_2_PhiReq/$entry
        Xexit_1724_symbol <= Xentry_1723_symbol; -- transition branch_block_stmt_134/bb_1_bb_2_PhiReq/$exit
        bb_1_bb_2_PhiReq_1722_symbol <= Xexit_1724_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_1_bb_2_PhiReq
      merge_stmt_180_PhiReqMerge_1725_symbol  <=  bb_1_bb_2_PhiReq_1722_symbol; -- place branch_block_stmt_134/merge_stmt_180_PhiReqMerge (optimized away) 
      merge_stmt_180_PhiAck_1726: Block -- branch_block_stmt_134/merge_stmt_180_PhiAck 
        signal merge_stmt_180_PhiAck_1726_start: Boolean;
        signal Xentry_1727_symbol: Boolean;
        signal Xexit_1728_symbol: Boolean;
        signal dummy_1729_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_180_PhiAck_1726_start <= merge_stmt_180_PhiReqMerge_1725_symbol; -- control passed to block
        Xentry_1727_symbol  <= merge_stmt_180_PhiAck_1726_start; -- transition branch_block_stmt_134/merge_stmt_180_PhiAck/$entry
        dummy_1729_symbol <= Xentry_1727_symbol; -- transition branch_block_stmt_134/merge_stmt_180_PhiAck/dummy
        Xexit_1728_symbol <= dummy_1729_symbol; -- transition branch_block_stmt_134/merge_stmt_180_PhiAck/$exit
        merge_stmt_180_PhiAck_1726_symbol <= Xexit_1728_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_180_PhiAck
      bb_1_bb_3_PhiReq_1730: Block -- branch_block_stmt_134/bb_1_bb_3_PhiReq 
        signal bb_1_bb_3_PhiReq_1730_start: Boolean;
        signal Xentry_1731_symbol: Boolean;
        signal Xexit_1732_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_3_PhiReq_1730_start <= bb_1_bb_3_552_symbol; -- control passed to block
        Xentry_1731_symbol  <= bb_1_bb_3_PhiReq_1730_start; -- transition branch_block_stmt_134/bb_1_bb_3_PhiReq/$entry
        Xexit_1732_symbol <= Xentry_1731_symbol; -- transition branch_block_stmt_134/bb_1_bb_3_PhiReq/$exit
        bb_1_bb_3_PhiReq_1730_symbol <= Xexit_1732_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_1_bb_3_PhiReq
      merge_stmt_227_PhiReqMerge_1733_symbol  <=  bb_1_bb_3_PhiReq_1730_symbol; -- place branch_block_stmt_134/merge_stmt_227_PhiReqMerge (optimized away) 
      merge_stmt_227_PhiAck_1734: Block -- branch_block_stmt_134/merge_stmt_227_PhiAck 
        signal merge_stmt_227_PhiAck_1734_start: Boolean;
        signal Xentry_1735_symbol: Boolean;
        signal Xexit_1736_symbol: Boolean;
        signal dummy_1737_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_227_PhiAck_1734_start <= merge_stmt_227_PhiReqMerge_1733_symbol; -- control passed to block
        Xentry_1735_symbol  <= merge_stmt_227_PhiAck_1734_start; -- transition branch_block_stmt_134/merge_stmt_227_PhiAck/$entry
        dummy_1737_symbol <= Xentry_1735_symbol; -- transition branch_block_stmt_134/merge_stmt_227_PhiAck/dummy
        Xexit_1736_symbol <= dummy_1737_symbol; -- transition branch_block_stmt_134/merge_stmt_227_PhiAck/$exit
        merge_stmt_227_PhiAck_1734_symbol <= Xexit_1736_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_227_PhiAck
      bb_3_bb_4_PhiReq_1738: Block -- branch_block_stmt_134/bb_3_bb_4_PhiReq 
        signal bb_3_bb_4_PhiReq_1738_start: Boolean;
        signal Xentry_1739_symbol: Boolean;
        signal Xexit_1740_symbol: Boolean;
        -- 
      begin -- 
        bb_3_bb_4_PhiReq_1738_start <= bb_3_bb_4_406_symbol; -- control passed to block
        Xentry_1739_symbol  <= bb_3_bb_4_PhiReq_1738_start; -- transition branch_block_stmt_134/bb_3_bb_4_PhiReq/$entry
        Xexit_1740_symbol <= Xentry_1739_symbol; -- transition branch_block_stmt_134/bb_3_bb_4_PhiReq/$exit
        bb_3_bb_4_PhiReq_1738_symbol <= Xexit_1740_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_3_bb_4_PhiReq
      bb_7_bb_4_PhiReq_1741: Block -- branch_block_stmt_134/bb_7_bb_4_PhiReq 
        signal bb_7_bb_4_PhiReq_1741_start: Boolean;
        signal Xentry_1742_symbol: Boolean;
        signal Xexit_1743_symbol: Boolean;
        -- 
      begin -- 
        bb_7_bb_4_PhiReq_1741_start <= bb_7_bb_4_432_symbol; -- control passed to block
        Xentry_1742_symbol  <= bb_7_bb_4_PhiReq_1741_start; -- transition branch_block_stmt_134/bb_7_bb_4_PhiReq/$entry
        Xexit_1743_symbol <= Xentry_1742_symbol; -- transition branch_block_stmt_134/bb_7_bb_4_PhiReq/$exit
        bb_7_bb_4_PhiReq_1741_symbol <= Xexit_1743_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_7_bb_4_PhiReq
      bb_8_bb_4_PhiReq_1744: Block -- branch_block_stmt_134/bb_8_bb_4_PhiReq 
        signal bb_8_bb_4_PhiReq_1744_start: Boolean;
        signal Xentry_1745_symbol: Boolean;
        signal Xexit_1746_symbol: Boolean;
        -- 
      begin -- 
        bb_8_bb_4_PhiReq_1744_start <= bb_8_bb_4_1446_symbol; -- control passed to block
        Xentry_1745_symbol  <= bb_8_bb_4_PhiReq_1744_start; -- transition branch_block_stmt_134/bb_8_bb_4_PhiReq/$entry
        Xexit_1746_symbol <= Xentry_1745_symbol; -- transition branch_block_stmt_134/bb_8_bb_4_PhiReq/$exit
        bb_8_bb_4_PhiReq_1744_symbol <= Xexit_1746_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_8_bb_4_PhiReq
      bb_9_bb_4_PhiReq_1747: Block -- branch_block_stmt_134/bb_9_bb_4_PhiReq 
        signal bb_9_bb_4_PhiReq_1747_start: Boolean;
        signal Xentry_1748_symbol: Boolean;
        signal Xexit_1749_symbol: Boolean;
        -- 
      begin -- 
        bb_9_bb_4_PhiReq_1747_start <= bb_9_bb_4_446_symbol; -- control passed to block
        Xentry_1748_symbol  <= bb_9_bb_4_PhiReq_1747_start; -- transition branch_block_stmt_134/bb_9_bb_4_PhiReq/$entry
        Xexit_1749_symbol <= Xentry_1748_symbol; -- transition branch_block_stmt_134/bb_9_bb_4_PhiReq/$exit
        bb_9_bb_4_PhiReq_1747_symbol <= Xexit_1749_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_9_bb_4_PhiReq
      merge_stmt_247_PhiReqMerge_1750_symbol  <=  bb_3_bb_4_PhiReq_1738_symbol or bb_7_bb_4_PhiReq_1741_symbol or bb_8_bb_4_PhiReq_1744_symbol or bb_9_bb_4_PhiReq_1747_symbol; -- place branch_block_stmt_134/merge_stmt_247_PhiReqMerge (optimized away) 
      merge_stmt_247_PhiAck_1751: Block -- branch_block_stmt_134/merge_stmt_247_PhiAck 
        signal merge_stmt_247_PhiAck_1751_start: Boolean;
        signal Xentry_1752_symbol: Boolean;
        signal Xexit_1753_symbol: Boolean;
        signal dummy_1754_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_247_PhiAck_1751_start <= merge_stmt_247_PhiReqMerge_1750_symbol; -- control passed to block
        Xentry_1752_symbol  <= merge_stmt_247_PhiAck_1751_start; -- transition branch_block_stmt_134/merge_stmt_247_PhiAck/$entry
        dummy_1754_symbol <= Xentry_1752_symbol; -- transition branch_block_stmt_134/merge_stmt_247_PhiAck/dummy
        Xexit_1753_symbol <= dummy_1754_symbol; -- transition branch_block_stmt_134/merge_stmt_247_PhiAck/$exit
        merge_stmt_247_PhiAck_1751_symbol <= Xexit_1753_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_247_PhiAck
      merge_stmt_280_dead_link_1755: Block -- branch_block_stmt_134/merge_stmt_280_dead_link 
        signal merge_stmt_280_dead_link_1755_start: Boolean;
        signal Xentry_1756_symbol: Boolean;
        signal Xexit_1757_symbol: Boolean;
        signal dead_transition_1758_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_280_dead_link_1755_start <= merge_stmt_280_x_xentry_x_xx_x416_symbol; -- control passed to block
        Xentry_1756_symbol  <= merge_stmt_280_dead_link_1755_start; -- transition branch_block_stmt_134/merge_stmt_280_dead_link/$entry
        dead_transition_1758_symbol <= false;
        Xexit_1757_symbol <= dead_transition_1758_symbol; -- transition branch_block_stmt_134/merge_stmt_280_dead_link/$exit
        merge_stmt_280_dead_link_1755_symbol <= Xexit_1757_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_280_dead_link
      bb_4_bb_5_PhiReq_1759: Block -- branch_block_stmt_134/bb_4_bb_5_PhiReq 
        signal bb_4_bb_5_PhiReq_1759_start: Boolean;
        signal Xentry_1760_symbol: Boolean;
        signal Xexit_1761_symbol: Boolean;
        -- 
      begin -- 
        bb_4_bb_5_PhiReq_1759_start <= bb_4_bb_5_1040_symbol; -- control passed to block
        Xentry_1760_symbol  <= bb_4_bb_5_PhiReq_1759_start; -- transition branch_block_stmt_134/bb_4_bb_5_PhiReq/$entry
        Xexit_1761_symbol <= Xentry_1760_symbol; -- transition branch_block_stmt_134/bb_4_bb_5_PhiReq/$exit
        bb_4_bb_5_PhiReq_1759_symbol <= Xexit_1761_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_4_bb_5_PhiReq
      merge_stmt_280_PhiReqMerge_1762_symbol  <=  bb_4_bb_5_PhiReq_1759_symbol; -- place branch_block_stmt_134/merge_stmt_280_PhiReqMerge (optimized away) 
      merge_stmt_280_PhiAck_1763: Block -- branch_block_stmt_134/merge_stmt_280_PhiAck 
        signal merge_stmt_280_PhiAck_1763_start: Boolean;
        signal Xentry_1764_symbol: Boolean;
        signal Xexit_1765_symbol: Boolean;
        signal dummy_1766_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_280_PhiAck_1763_start <= merge_stmt_280_PhiReqMerge_1762_symbol; -- control passed to block
        Xentry_1764_symbol  <= merge_stmt_280_PhiAck_1763_start; -- transition branch_block_stmt_134/merge_stmt_280_PhiAck/$entry
        dummy_1766_symbol <= Xentry_1764_symbol; -- transition branch_block_stmt_134/merge_stmt_280_PhiAck/dummy
        Xexit_1765_symbol <= dummy_1766_symbol; -- transition branch_block_stmt_134/merge_stmt_280_PhiAck/$exit
        merge_stmt_280_PhiAck_1763_symbol <= Xexit_1765_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_280_PhiAck
      merge_stmt_304_dead_link_1767: Block -- branch_block_stmt_134/merge_stmt_304_dead_link 
        signal merge_stmt_304_dead_link_1767_start: Boolean;
        signal Xentry_1768_symbol: Boolean;
        signal Xexit_1769_symbol: Boolean;
        signal dead_transition_1770_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_304_dead_link_1767_start <= merge_stmt_304_x_xentry_x_xx_x422_symbol; -- control passed to block
        Xentry_1768_symbol  <= merge_stmt_304_dead_link_1767_start; -- transition branch_block_stmt_134/merge_stmt_304_dead_link/$entry
        dead_transition_1770_symbol <= false;
        Xexit_1769_symbol <= dead_transition_1770_symbol; -- transition branch_block_stmt_134/merge_stmt_304_dead_link/$exit
        merge_stmt_304_dead_link_1767_symbol <= Xexit_1769_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_304_dead_link
      bb_5_bb_6_PhiReq_1771: Block -- branch_block_stmt_134/bb_5_bb_6_PhiReq 
        signal bb_5_bb_6_PhiReq_1771_start: Boolean;
        signal Xentry_1772_symbol: Boolean;
        signal Xexit_1773_symbol: Boolean;
        -- 
      begin -- 
        bb_5_bb_6_PhiReq_1771_start <= bb_5_bb_6_1173_symbol; -- control passed to block
        Xentry_1772_symbol  <= bb_5_bb_6_PhiReq_1771_start; -- transition branch_block_stmt_134/bb_5_bb_6_PhiReq/$entry
        Xexit_1773_symbol <= Xentry_1772_symbol; -- transition branch_block_stmt_134/bb_5_bb_6_PhiReq/$exit
        bb_5_bb_6_PhiReq_1771_symbol <= Xexit_1773_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_5_bb_6_PhiReq
      merge_stmt_304_PhiReqMerge_1774_symbol  <=  bb_5_bb_6_PhiReq_1771_symbol; -- place branch_block_stmt_134/merge_stmt_304_PhiReqMerge (optimized away) 
      merge_stmt_304_PhiAck_1775: Block -- branch_block_stmt_134/merge_stmt_304_PhiAck 
        signal merge_stmt_304_PhiAck_1775_start: Boolean;
        signal Xentry_1776_symbol: Boolean;
        signal Xexit_1777_symbol: Boolean;
        signal dummy_1778_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_304_PhiAck_1775_start <= merge_stmt_304_PhiReqMerge_1774_symbol; -- control passed to block
        Xentry_1776_symbol  <= merge_stmt_304_PhiAck_1775_start; -- transition branch_block_stmt_134/merge_stmt_304_PhiAck/$entry
        dummy_1778_symbol <= Xentry_1776_symbol; -- transition branch_block_stmt_134/merge_stmt_304_PhiAck/dummy
        Xexit_1777_symbol <= dummy_1778_symbol; -- transition branch_block_stmt_134/merge_stmt_304_PhiAck/$exit
        merge_stmt_304_PhiAck_1775_symbol <= Xexit_1777_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_304_PhiAck
      bb_5_bb_7_PhiReq_1779: Block -- branch_block_stmt_134/bb_5_bb_7_PhiReq 
        signal bb_5_bb_7_PhiReq_1779_start: Boolean;
        signal Xentry_1780_symbol: Boolean;
        signal Xexit_1781_symbol: Boolean;
        -- 
      begin -- 
        bb_5_bb_7_PhiReq_1779_start <= bb_5_bb_7_1174_symbol; -- control passed to block
        Xentry_1780_symbol  <= bb_5_bb_7_PhiReq_1779_start; -- transition branch_block_stmt_134/bb_5_bb_7_PhiReq/$entry
        Xexit_1781_symbol <= Xentry_1780_symbol; -- transition branch_block_stmt_134/bb_5_bb_7_PhiReq/$exit
        bb_5_bb_7_PhiReq_1779_symbol <= Xexit_1781_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_5_bb_7_PhiReq
      bb_6_bb_7_PhiReq_1782: Block -- branch_block_stmt_134/bb_6_bb_7_PhiReq 
        signal bb_6_bb_7_PhiReq_1782_start: Boolean;
        signal Xentry_1783_symbol: Boolean;
        signal Xexit_1784_symbol: Boolean;
        -- 
      begin -- 
        bb_6_bb_7_PhiReq_1782_start <= bb_6_bb_7_426_symbol; -- control passed to block
        Xentry_1783_symbol  <= bb_6_bb_7_PhiReq_1782_start; -- transition branch_block_stmt_134/bb_6_bb_7_PhiReq/$entry
        Xexit_1784_symbol <= Xentry_1783_symbol; -- transition branch_block_stmt_134/bb_6_bb_7_PhiReq/$exit
        bb_6_bb_7_PhiReq_1782_symbol <= Xexit_1784_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_6_bb_7_PhiReq
      merge_stmt_321_PhiReqMerge_1785_symbol  <=  bb_5_bb_7_PhiReq_1779_symbol or bb_6_bb_7_PhiReq_1782_symbol; -- place branch_block_stmt_134/merge_stmt_321_PhiReqMerge (optimized away) 
      merge_stmt_321_PhiAck_1786: Block -- branch_block_stmt_134/merge_stmt_321_PhiAck 
        signal merge_stmt_321_PhiAck_1786_start: Boolean;
        signal Xentry_1787_symbol: Boolean;
        signal Xexit_1788_symbol: Boolean;
        signal dummy_1789_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_321_PhiAck_1786_start <= merge_stmt_321_PhiReqMerge_1785_symbol; -- control passed to block
        Xentry_1787_symbol  <= merge_stmt_321_PhiAck_1786_start; -- transition branch_block_stmt_134/merge_stmt_321_PhiAck/$entry
        dummy_1789_symbol <= Xentry_1787_symbol; -- transition branch_block_stmt_134/merge_stmt_321_PhiAck/dummy
        Xexit_1788_symbol <= dummy_1789_symbol; -- transition branch_block_stmt_134/merge_stmt_321_PhiAck/$exit
        merge_stmt_321_PhiAck_1786_symbol <= Xexit_1788_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_321_PhiAck
      bb_4_bb_8_PhiReq_1790: Block -- branch_block_stmt_134/bb_4_bb_8_PhiReq 
        signal bb_4_bb_8_PhiReq_1790_start: Boolean;
        signal Xentry_1791_symbol: Boolean;
        signal Xexit_1792_symbol: Boolean;
        -- 
      begin -- 
        bb_4_bb_8_PhiReq_1790_start <= bb_4_bb_8_1041_symbol; -- control passed to block
        Xentry_1791_symbol  <= bb_4_bb_8_PhiReq_1790_start; -- transition branch_block_stmt_134/bb_4_bb_8_PhiReq/$entry
        Xexit_1792_symbol <= Xentry_1791_symbol; -- transition branch_block_stmt_134/bb_4_bb_8_PhiReq/$exit
        bb_4_bb_8_PhiReq_1790_symbol <= Xexit_1792_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_4_bb_8_PhiReq
      merge_stmt_340_PhiReqMerge_1793_symbol  <=  bb_4_bb_8_PhiReq_1790_symbol; -- place branch_block_stmt_134/merge_stmt_340_PhiReqMerge (optimized away) 
      merge_stmt_340_PhiAck_1794: Block -- branch_block_stmt_134/merge_stmt_340_PhiAck 
        signal merge_stmt_340_PhiAck_1794_start: Boolean;
        signal Xentry_1795_symbol: Boolean;
        signal Xexit_1796_symbol: Boolean;
        signal dummy_1797_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_340_PhiAck_1794_start <= merge_stmt_340_PhiReqMerge_1793_symbol; -- control passed to block
        Xentry_1795_symbol  <= merge_stmt_340_PhiAck_1794_start; -- transition branch_block_stmt_134/merge_stmt_340_PhiAck/$entry
        dummy_1797_symbol <= Xentry_1795_symbol; -- transition branch_block_stmt_134/merge_stmt_340_PhiAck/dummy
        Xexit_1796_symbol <= dummy_1797_symbol; -- transition branch_block_stmt_134/merge_stmt_340_PhiAck/$exit
        merge_stmt_340_PhiAck_1794_symbol <= Xexit_1796_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_340_PhiAck
      merge_stmt_360_dead_link_1798: Block -- branch_block_stmt_134/merge_stmt_360_dead_link 
        signal merge_stmt_360_dead_link_1798_start: Boolean;
        signal Xentry_1799_symbol: Boolean;
        signal Xexit_1800_symbol: Boolean;
        signal dead_transition_1801_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_360_dead_link_1798_start <= merge_stmt_360_x_xentry_x_xx_x438_symbol; -- control passed to block
        Xentry_1799_symbol  <= merge_stmt_360_dead_link_1798_start; -- transition branch_block_stmt_134/merge_stmt_360_dead_link/$entry
        dead_transition_1801_symbol <= false;
        Xexit_1800_symbol <= dead_transition_1801_symbol; -- transition branch_block_stmt_134/merge_stmt_360_dead_link/$exit
        merge_stmt_360_dead_link_1798_symbol <= Xexit_1800_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_360_dead_link
      bb_8_bb_9_PhiReq_1802: Block -- branch_block_stmt_134/bb_8_bb_9_PhiReq 
        signal bb_8_bb_9_PhiReq_1802_start: Boolean;
        signal Xentry_1803_symbol: Boolean;
        signal Xexit_1804_symbol: Boolean;
        -- 
      begin -- 
        bb_8_bb_9_PhiReq_1802_start <= bb_8_bb_9_1445_symbol; -- control passed to block
        Xentry_1803_symbol  <= bb_8_bb_9_PhiReq_1802_start; -- transition branch_block_stmt_134/bb_8_bb_9_PhiReq/$entry
        Xexit_1804_symbol <= Xentry_1803_symbol; -- transition branch_block_stmt_134/bb_8_bb_9_PhiReq/$exit
        bb_8_bb_9_PhiReq_1802_symbol <= Xexit_1804_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/bb_8_bb_9_PhiReq
      merge_stmt_360_PhiReqMerge_1805_symbol  <=  bb_8_bb_9_PhiReq_1802_symbol; -- place branch_block_stmt_134/merge_stmt_360_PhiReqMerge (optimized away) 
      merge_stmt_360_PhiAck_1806: Block -- branch_block_stmt_134/merge_stmt_360_PhiAck 
        signal merge_stmt_360_PhiAck_1806_start: Boolean;
        signal Xentry_1807_symbol: Boolean;
        signal Xexit_1808_symbol: Boolean;
        signal dummy_1809_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_360_PhiAck_1806_start <= merge_stmt_360_PhiReqMerge_1805_symbol; -- control passed to block
        Xentry_1807_symbol  <= merge_stmt_360_PhiAck_1806_start; -- transition branch_block_stmt_134/merge_stmt_360_PhiAck/$entry
        dummy_1809_symbol <= Xentry_1807_symbol; -- transition branch_block_stmt_134/merge_stmt_360_PhiAck/dummy
        Xexit_1808_symbol <= dummy_1809_symbol; -- transition branch_block_stmt_134/merge_stmt_360_PhiAck/$exit
        merge_stmt_360_PhiAck_1806_symbol <= Xexit_1808_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_134/merge_stmt_360_PhiAck
      Xexit_387_symbol <= branch_block_stmt_134_x_xexit_x_xx_x389_symbol; -- transition branch_block_stmt_134/$exit
      branch_block_stmt_134_385_symbol <= Xexit_387_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_134
    Xexit_384_symbol <= branch_block_stmt_134_385_symbol; -- transition $exit
    fin  <=  '1' when Xexit_384_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_192_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_192_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_192_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_192_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_201_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_201_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_201_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_201_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_207_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_207_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_311_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_311_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_388_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_388_root_address : std_logic_vector(2 downto 0);
    signal command_146 : std_logic_vector(31 downto 0);
    signal expr_157_wire_constant : std_logic_vector(31 downto 0);
    signal expr_187_wire_constant : std_logic_vector(31 downto 0);
    signal expr_219_wire_constant : std_logic_vector(31 downto 0);
    signal expr_236_wire_constant : std_logic_vector(31 downto 0);
    signal expr_271_wire_constant : std_logic_vector(31 downto 0);
    signal expr_351_wire_constant : std_logic_vector(31 downto 0);
    signal iNsTr_10_208 : std_logic_vector(31 downto 0);
    signal iNsTr_12_216 : std_logic_vector(31 downto 0);
    signal iNsTr_13_221 : std_logic_vector(31 downto 0);
    signal iNsTr_16_233 : std_logic_vector(31 downto 0);
    signal iNsTr_18_242 : std_logic_vector(31 downto 0);
    signal iNsTr_21_252 : std_logic_vector(31 downto 0);
    signal iNsTr_22_256 : std_logic_vector(7 downto 0);
    signal iNsTr_24_264 : std_logic_vector(7 downto 0);
    signal iNsTr_25_268 : std_logic_vector(31 downto 0);
    signal iNsTr_26_273 : std_logic_vector(0 downto 0);
    signal iNsTr_28_283 : std_logic_vector(31 downto 0);
    signal iNsTr_2_164 : std_logic_vector(31 downto 0);
    signal iNsTr_30_290 : std_logic_vector(31 downto 0);
    signal iNsTr_31_297 : std_logic_vector(0 downto 0);
    signal iNsTr_33_344 : std_logic_vector(7 downto 0);
    signal iNsTr_34_348 : std_logic_vector(31 downto 0);
    signal iNsTr_35_353 : std_logic_vector(0 downto 0);
    signal iNsTr_37_307 : std_logic_vector(31 downto 0);
    signal iNsTr_38_312 : std_logic_vector(31 downto 0);
    signal iNsTr_39_316 : std_logic_vector(31 downto 0);
    signal iNsTr_3_173 : std_logic_vector(0 downto 0);
    signal iNsTr_42_325 : std_logic_vector(31 downto 0);
    signal iNsTr_43_329 : std_logic_vector(31 downto 0);
    signal iNsTr_44_334 : std_logic_vector(31 downto 0);
    signal iNsTr_47_365 : std_logic_vector(31 downto 0);
    signal iNsTr_48_369 : std_logic_vector(31 downto 0);
    signal iNsTr_49_373 : std_logic_vector(31 downto 0);
    signal iNsTr_51_380 : std_logic_vector(31 downto 0);
    signal iNsTr_52_384 : std_logic_vector(31 downto 0);
    signal iNsTr_53_389 : std_logic_vector(31 downto 0);
    signal iNsTr_55_397 : std_logic_vector(31 downto 0);
    signal iNsTr_5_184 : std_logic_vector(31 downto 0);
    signal iNsTr_6_189 : std_logic_vector(31 downto 0);
    signal iNsTr_7_194 : std_logic_vector(31 downto 0);
    signal iNsTr_8_198 : std_logic_vector(31 downto 0);
    signal iNsTr_9_203 : std_logic_vector(31 downto 0);
    signal i_142 : std_logic_vector(31 downto 0);
    signal ptr_deref_156_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_156_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_156_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_163_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_163_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_183_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_183_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_197_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_197_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_210_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_210_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_210_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_210_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_210_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_210_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_215_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_215_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_223_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_223_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_223_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_235_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_235_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_235_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_258_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_258_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_258_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_263_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_263_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_285_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_285_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_285_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_315_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_315_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_315_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_315_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_315_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_324_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_324_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_343_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_343_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_375_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_375_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_375_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_383_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_383_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_391_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_391_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_391_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_391_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_391_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_391_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_396_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_396_word_address_0 : std_logic_vector(0 downto 0);
    signal put_link_154 : std_logic_vector(31 downto 0);
    signal ret_150 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_191_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_191_scaled : std_logic_vector(2 downto 0);
    signal simple_obj_ref_200_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_200_scaled : std_logic_vector(2 downto 0);
    signal simple_obj_ref_243_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_243_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_254_wire : std_logic_vector(7 downto 0);
    signal simple_obj_ref_282_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_282_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_289_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_289_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_306_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_306_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_317_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_317_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_367_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_379_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_379_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_398_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_398_word_address_0 : std_logic_vector(0 downto 0);
    signal type_cast_168_wire : std_logic_vector(31 downto 0);
    signal type_cast_170_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_293_wire : std_logic_vector(31 downto 0);
    signal type_cast_295_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_337_wire : std_logic_vector(31 downto 0);
    signal xxfree_queue_managerxxbodyxxcommand_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxfree_queue_managerxxbodyxxi_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxfree_queue_managerxxbodyxxput_link_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxfree_queue_managerxxbodyxxret_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_192_offset_scale_factor_0 <= "010";
    array_obj_ref_192_resized_base_address <= "000";
    array_obj_ref_201_offset_scale_factor_0 <= "010";
    array_obj_ref_201_resized_base_address <= "000";
    command_146 <= "00000000000000000000000000000000";
    expr_157_wire_constant <= "00000000000000000000000000000000";
    expr_187_wire_constant <= "00000000000000000000000000000001";
    expr_219_wire_constant <= "00000000000000000000000000000001";
    expr_236_wire_constant <= "11111111111111111111111111111111";
    expr_271_wire_constant <= "00000000000000000000000000000010";
    expr_351_wire_constant <= "00000000000000000000000000000001";
    iNsTr_16_233 <= "00000000000000000000000000000010";
    iNsTr_18_242 <= "00000000000000000000000000000000";
    iNsTr_21_252 <= "00000000000000000000000000000000";
    iNsTr_44_334 <= "00000000000000000000000000000000";
    iNsTr_47_365 <= "00000000000000000000000000000000";
    i_142 <= "00000000000000000000000000000000";
    ptr_deref_156_word_address_0 <= "0";
    ptr_deref_163_word_address_0 <= "0";
    ptr_deref_183_word_address_0 <= "0";
    ptr_deref_197_word_address_0 <= "0";
    ptr_deref_210_word_offset_0 <= "000";
    ptr_deref_215_word_address_0 <= "0";
    ptr_deref_223_word_address_0 <= "0";
    ptr_deref_235_word_address_0 <= "010";
    ptr_deref_258_word_address_0 <= "0";
    ptr_deref_263_word_address_0 <= "0";
    ptr_deref_285_word_address_0 <= "0";
    ptr_deref_315_word_offset_0 <= "000";
    ptr_deref_324_word_address_0 <= "0";
    ptr_deref_343_word_address_0 <= "0";
    ptr_deref_375_word_address_0 <= "0";
    ptr_deref_383_word_address_0 <= "0";
    ptr_deref_391_word_offset_0 <= "000";
    ptr_deref_396_word_address_0 <= "0";
    put_link_154 <= "00000000000000000000000000000000";
    ret_150 <= "00000000000000000000000000000000";
    simple_obj_ref_243_word_address_0 <= "0";
    simple_obj_ref_282_word_address_0 <= "0";
    simple_obj_ref_289_word_address_0 <= "0";
    simple_obj_ref_306_word_address_0 <= "0";
    simple_obj_ref_317_word_address_0 <= "0";
    simple_obj_ref_379_word_address_0 <= "0";
    simple_obj_ref_398_word_address_0 <= "0";
    type_cast_170_wire_constant <= "00000000000000000000000000000001";
    type_cast_295_wire_constant <= "11111111111111111111111111111111";
    xxfree_queue_managerxxbodyxxcommand_alloc_base_address <= "0";
    xxfree_queue_managerxxbodyxxi_alloc_base_address <= "0";
    xxfree_queue_managerxxbodyxxput_link_alloc_base_address <= "0";
    xxfree_queue_managerxxbodyxxret_alloc_base_address <= "0";
    addr_of_193_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_192_root_address, dout => iNsTr_7_194, req => addr_of_193_final_reg_req_0, ack => addr_of_193_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_202_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_201_root_address, dout => iNsTr_9_203, req => addr_of_202_final_reg_req_0, ack => addr_of_202_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_192_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_6_189, dout => simple_obj_ref_191_resized, req => array_obj_ref_192_index_0_resize_req_0, ack => array_obj_ref_192_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_192_offset_inst: RegisterBase generic map(in_data_width => 3,out_data_width => 3) -- 
      port map( din => simple_obj_ref_191_scaled, dout => array_obj_ref_192_final_offset, req => array_obj_ref_192_offset_inst_req_0, ack => array_obj_ref_192_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_201_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_8_198, dout => simple_obj_ref_200_resized, req => array_obj_ref_201_index_0_resize_req_0, ack => array_obj_ref_201_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_201_offset_inst: RegisterBase generic map(in_data_width => 3,out_data_width => 3) -- 
      port map( din => simple_obj_ref_200_scaled, dout => array_obj_ref_201_final_offset, req => array_obj_ref_201_offset_inst_req_0, ack => array_obj_ref_201_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_207_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_9_203, dout => array_obj_ref_207_resized_base_address, req => array_obj_ref_207_base_resize_req_0, ack => array_obj_ref_207_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_207_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_207_root_address, dout => iNsTr_10_208, req => array_obj_ref_207_final_reg_req_0, ack => array_obj_ref_207_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_311_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_37_307, dout => array_obj_ref_311_resized_base_address, req => array_obj_ref_311_base_resize_req_0, ack => array_obj_ref_311_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_311_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_311_root_address, dout => iNsTr_38_312, req => array_obj_ref_311_final_reg_req_0, ack => array_obj_ref_311_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_388_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_52_384, dout => array_obj_ref_388_resized_base_address, req => array_obj_ref_388_base_resize_req_0, ack => array_obj_ref_388_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_388_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_388_root_address, dout => iNsTr_53_389, req => array_obj_ref_388_final_reg_req_0, ack => array_obj_ref_388_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_210_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_10_208, dout => ptr_deref_210_resized_base_address, req => ptr_deref_210_base_resize_req_0, ack => ptr_deref_210_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_315_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_38_312, dout => ptr_deref_315_resized_base_address, req => ptr_deref_315_base_resize_req_0, ack => ptr_deref_315_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_391_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_53_389, dout => ptr_deref_391_resized_base_address, req => ptr_deref_391_base_resize_req_0, ack => ptr_deref_391_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_168_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_2_164, dout => type_cast_168_wire, req => type_cast_168_inst_req_0, ack => type_cast_168_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_255_inst: RegisterBase generic map(in_data_width => 8,out_data_width => 8) -- 
      port map( din => simple_obj_ref_254_wire, dout => iNsTr_22_256, req => type_cast_255_inst_req_0, ack => type_cast_255_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_267_inst: RegisterBase generic map(in_data_width => 8,out_data_width => 32) -- 
      port map( din => iNsTr_24_264, dout => iNsTr_25_268, req => type_cast_267_inst_req_0, ack => type_cast_267_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_293_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_30_290, dout => type_cast_293_wire, req => type_cast_293_inst_req_0, ack => type_cast_293_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_328_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_42_325, dout => iNsTr_43_329, req => type_cast_328_inst_req_0, ack => type_cast_328_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_337_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_43_329, dout => type_cast_337_wire, req => type_cast_337_inst_req_0, ack => type_cast_337_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_347_inst: RegisterBase generic map(in_data_width => 8,out_data_width => 32) -- 
      port map( din => iNsTr_33_344, dout => iNsTr_34_348, req => type_cast_347_inst_req_0, ack => type_cast_347_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_368_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_367_wire, dout => iNsTr_48_369, req => type_cast_368_inst_req_0, ack => type_cast_368_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_372_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_48_369, dout => iNsTr_49_373, req => type_cast_372_inst_req_0, ack => type_cast_372_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_192_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_192_root_address_inst_ack_0 <= array_obj_ref_192_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_192_final_offset;
      array_obj_ref_192_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_201_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_201_root_address_inst_ack_0 <= array_obj_ref_201_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_201_final_offset;
      array_obj_ref_201_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_207_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_207_root_address_inst_ack_0 <= array_obj_ref_207_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_207_resized_base_address;
      array_obj_ref_207_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_311_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_311_root_address_inst_ack_0 <= array_obj_ref_311_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_311_resized_base_address;
      array_obj_ref_311_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_388_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_388_root_address_inst_ack_0 <= array_obj_ref_388_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_388_resized_base_address;
      array_obj_ref_388_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_156_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_156_gather_scatter_ack_0 <= ptr_deref_156_gather_scatter_req_0;
      aggregated_sig <= expr_157_wire_constant;
      ptr_deref_156_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_163_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_163_gather_scatter_ack_0 <= ptr_deref_163_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_163_data_0;
      iNsTr_2_164 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_183_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_183_gather_scatter_ack_0 <= ptr_deref_183_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_183_data_0;
      iNsTr_5_184 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_197_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_197_gather_scatter_ack_0 <= ptr_deref_197_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_197_data_0;
      iNsTr_8_198 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_210_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_210_addr_0_ack_0 <= ptr_deref_210_addr_0_req_0;
      aggregated_sig <= ptr_deref_210_root_address;
      ptr_deref_210_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_210_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_210_gather_scatter_ack_0 <= ptr_deref_210_gather_scatter_req_0;
      aggregated_sig <= iNsTr_7_194;
      ptr_deref_210_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_210_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_210_root_address_inst_ack_0 <= ptr_deref_210_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_210_resized_base_address;
      ptr_deref_210_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_215_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_215_gather_scatter_ack_0 <= ptr_deref_215_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_215_data_0;
      iNsTr_12_216 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_223_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_223_gather_scatter_ack_0 <= ptr_deref_223_gather_scatter_req_0;
      aggregated_sig <= iNsTr_13_221;
      ptr_deref_223_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_235_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_235_gather_scatter_ack_0 <= ptr_deref_235_gather_scatter_req_0;
      aggregated_sig <= expr_236_wire_constant;
      ptr_deref_235_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_258_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_258_gather_scatter_ack_0 <= ptr_deref_258_gather_scatter_req_0;
      aggregated_sig <= iNsTr_22_256;
      ptr_deref_258_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_263_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_263_gather_scatter_ack_0 <= ptr_deref_263_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_263_data_0;
      iNsTr_24_264 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_285_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_285_gather_scatter_ack_0 <= ptr_deref_285_gather_scatter_req_0;
      aggregated_sig <= iNsTr_28_283;
      ptr_deref_285_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_315_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_315_addr_0_ack_0 <= ptr_deref_315_addr_0_req_0;
      aggregated_sig <= ptr_deref_315_root_address;
      ptr_deref_315_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_315_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_315_gather_scatter_ack_0 <= ptr_deref_315_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_315_data_0;
      iNsTr_39_316 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_315_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_315_root_address_inst_ack_0 <= ptr_deref_315_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_315_resized_base_address;
      ptr_deref_315_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_324_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_324_gather_scatter_ack_0 <= ptr_deref_324_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_324_data_0;
      iNsTr_42_325 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_343_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_343_gather_scatter_ack_0 <= ptr_deref_343_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_343_data_0;
      iNsTr_33_344 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_375_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_375_gather_scatter_ack_0 <= ptr_deref_375_gather_scatter_req_0;
      aggregated_sig <= iNsTr_49_373;
      ptr_deref_375_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_383_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_383_gather_scatter_ack_0 <= ptr_deref_383_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_383_data_0;
      iNsTr_52_384 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_391_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_391_addr_0_ack_0 <= ptr_deref_391_addr_0_req_0;
      aggregated_sig <= ptr_deref_391_root_address;
      ptr_deref_391_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_391_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_391_gather_scatter_ack_0 <= ptr_deref_391_gather_scatter_req_0;
      aggregated_sig <= iNsTr_51_380;
      ptr_deref_391_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_391_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_391_root_address_inst_ack_0 <= ptr_deref_391_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_391_resized_base_address;
      ptr_deref_391_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_396_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_396_gather_scatter_ack_0 <= ptr_deref_396_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_396_data_0;
      iNsTr_55_397 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_243_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_243_gather_scatter_ack_0 <= simple_obj_ref_243_gather_scatter_req_0;
      aggregated_sig <= iNsTr_18_242;
      simple_obj_ref_243_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_282_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_282_gather_scatter_ack_0 <= simple_obj_ref_282_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_282_data_0;
      iNsTr_28_283 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_289_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_289_gather_scatter_ack_0 <= simple_obj_ref_289_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_289_data_0;
      iNsTr_30_290 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_306_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_306_gather_scatter_ack_0 <= simple_obj_ref_306_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_306_data_0;
      iNsTr_37_307 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_317_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_317_gather_scatter_ack_0 <= simple_obj_ref_317_gather_scatter_req_0;
      aggregated_sig <= iNsTr_39_316;
      simple_obj_ref_317_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_379_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_379_gather_scatter_ack_0 <= simple_obj_ref_379_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_379_data_0;
      iNsTr_51_380 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_398_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_398_gather_scatter_ack_0 <= simple_obj_ref_398_gather_scatter_req_0;
      aggregated_sig <= iNsTr_55_397;
      simple_obj_ref_398_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_174_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_3_173;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_174_branch_req_0,
          ack0 => if_stmt_174_branch_ack_0,
          ack1 => if_stmt_174_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_274_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_26_273;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_274_branch_req_0,
          ack0 => if_stmt_274_branch_ack_0,
          ack1 => if_stmt_274_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_298_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_31_297;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_298_branch_req_0,
          ack0 => if_stmt_298_branch_ack_0,
          ack1 => if_stmt_298_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_354_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_35_353;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_354_branch_req_0,
          ack0 => if_stmt_354_branch_ack_0,
          ack1 => if_stmt_354_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_192_index_0_scale 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_191_resized;
      simple_obj_ref_191_scaled <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_192_index_0_scale_req_0,
          ackL => array_obj_ref_192_index_0_scale_ack_0,
          reqR => array_obj_ref_192_index_0_scale_req_1,
          ackR => array_obj_ref_192_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_201_index_0_scale 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_200_resized;
      simple_obj_ref_200_scaled <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_201_index_0_scale_req_0,
          ackL => array_obj_ref_201_index_0_scale_ack_0,
          reqR => array_obj_ref_201_index_0_scale_req_1,
          ackR => array_obj_ref_201_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_171_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_168_wire;
      iNsTr_3_173 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_171_inst_req_0,
          ackL => binary_171_inst_ack_0,
          reqR => binary_171_inst_req_1,
          ackR => binary_171_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_188_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_5_184;
      iNsTr_6_189 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_188_inst_req_0,
          ackL => binary_188_inst_ack_0,
          reqR => binary_188_inst_req_1,
          ackR => binary_188_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_220_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_12_216;
      iNsTr_13_221 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_220_inst_req_0,
          ackL => binary_220_inst_ack_0,
          reqR => binary_220_inst_req_1,
          ackR => binary_220_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_272_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_25_268;
      iNsTr_26_273 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000010",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_272_inst_req_0,
          ackL => binary_272_inst_ack_0,
          reqR => binary_272_inst_req_1,
          ackR => binary_272_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_296_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_293_wire;
      iNsTr_31_297 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_296_inst_req_0,
          ackL => binary_296_inst_ack_0,
          reqR => binary_296_inst_req_1,
          ackR => binary_296_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_352_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_34_348;
      iNsTr_35_353 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_352_inst_req_0,
          ackL => binary_352_inst_ack_0,
          reqR => binary_352_inst_req_1,
          ackR => binary_352_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared load operator group (0) : ptr_deref_163_load_0 ptr_deref_183_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_163_load_0_req_0;
      reqL(0) <= ptr_deref_183_load_0_req_0;
      ptr_deref_163_load_0_ack_0 <= ackL(1);
      ptr_deref_183_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_163_load_0_req_1;
      reqR(0) <= ptr_deref_183_load_0_req_1;
      ptr_deref_163_load_0_ack_1 <= ackR(1);
      ptr_deref_183_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_163_word_address_0 & ptr_deref_183_word_address_0;
      ptr_deref_163_data_0 <= data_out(63 downto 32);
      ptr_deref_183_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_11_lr_req(2),
          mack => memory_space_11_lr_ack(2),
          maddr => memory_space_11_lr_addr(2 downto 2),
          mtag => memory_space_11_lr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_11_lc_req(2),
          mack => memory_space_11_lc_ack(2),
          mdata => memory_space_11_lc_data(95 downto 64),
          mtag => memory_space_11_lc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_197_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_197_load_0_req_0;
      ptr_deref_197_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_197_load_0_req_1;
      ptr_deref_197_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_197_word_address_0;
      ptr_deref_197_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_11_lr_req(1),
          mack => memory_space_11_lr_ack(1),
          maddr => memory_space_11_lr_addr(1 downto 1),
          mtag => memory_space_11_lr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_11_lc_req(1),
          mack => memory_space_11_lc_ack(1),
          mdata => memory_space_11_lc_data(63 downto 32),
          mtag => memory_space_11_lc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_215_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_215_load_0_req_0;
      ptr_deref_215_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_215_load_0_req_1;
      ptr_deref_215_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_215_word_address_0;
      ptr_deref_215_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_11_lr_req(0),
          mack => memory_space_11_lr_ack(0),
          maddr => memory_space_11_lr_addr(0 downto 0),
          mtag => memory_space_11_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_11_lc_req(0),
          mack => memory_space_11_lc_ack(0),
          mdata => memory_space_11_lc_data(31 downto 0),
          mtag => memory_space_11_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_263_load_0 ptr_deref_343_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_263_load_0_req_0;
      reqL(0) <= ptr_deref_343_load_0_req_0;
      ptr_deref_263_load_0_ack_0 <= ackL(1);
      ptr_deref_343_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_263_load_0_req_1;
      reqR(0) <= ptr_deref_343_load_0_req_1;
      ptr_deref_263_load_0_ack_1 <= ackR(1);
      ptr_deref_343_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_263_word_address_0 & ptr_deref_343_word_address_0;
      ptr_deref_263_data_0 <= data_out(15 downto 8);
      ptr_deref_343_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_12_lr_req(0),
          mack => memory_space_12_lr_ack(0),
          maddr => memory_space_12_lr_addr(0 downto 0),
          mtag => memory_space_12_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_12_lc_req(0),
          mack => memory_space_12_lc_ack(0),
          mdata => memory_space_12_lc_data(7 downto 0),
          mtag => memory_space_12_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_315_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_315_load_0_req_0;
      ptr_deref_315_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_315_load_0_req_1;
      ptr_deref_315_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_315_word_address_0;
      ptr_deref_315_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 3,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(2 downto 0),
          mtag => memory_space_1_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_324_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_324_load_0_req_0;
      ptr_deref_324_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_324_load_0_req_1;
      ptr_deref_324_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_324_word_address_0;
      ptr_deref_324_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_13_lr_req(0),
          mack => memory_space_13_lr_ack(0),
          maddr => memory_space_13_lr_addr(0 downto 0),
          mtag => memory_space_13_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_13_lc_req(0),
          mack => memory_space_13_lc_ack(0),
          mdata => memory_space_13_lc_data(31 downto 0),
          mtag => memory_space_13_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_383_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_383_load_0_req_0;
      ptr_deref_383_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_383_load_0_req_1;
      ptr_deref_383_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_383_word_address_0;
      ptr_deref_383_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_14_lr_req(1),
          mack => memory_space_14_lr_ack(1),
          maddr => memory_space_14_lr_addr(1 downto 1),
          mtag => memory_space_14_lr_tag(1 downto 1),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_14_lc_req(1),
          mack => memory_space_14_lc_ack(1),
          mdata => memory_space_14_lc_data(63 downto 32),
          mtag => memory_space_14_lc_tag(1 downto 1),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_396_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_396_load_0_req_0;
      ptr_deref_396_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_396_load_0_req_1;
      ptr_deref_396_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_396_word_address_0;
      ptr_deref_396_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_14_lr_req(0),
          mack => memory_space_14_lr_ack(0),
          maddr => memory_space_14_lr_addr(0 downto 0),
          mtag => memory_space_14_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_14_lc_req(0),
          mack => memory_space_14_lc_ack(0),
          mdata => memory_space_14_lc_data(31 downto 0),
          mtag => memory_space_14_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared load operator group (8) : simple_obj_ref_379_load_0 simple_obj_ref_282_load_0 simple_obj_ref_306_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= simple_obj_ref_379_load_0_req_0;
      reqL(1) <= simple_obj_ref_282_load_0_req_0;
      reqL(0) <= simple_obj_ref_306_load_0_req_0;
      simple_obj_ref_379_load_0_ack_0 <= ackL(2);
      simple_obj_ref_282_load_0_ack_0 <= ackL(1);
      simple_obj_ref_306_load_0_ack_0 <= ackL(0);
      reqR(2) <= simple_obj_ref_379_load_0_req_1;
      reqR(1) <= simple_obj_ref_282_load_0_req_1;
      reqR(0) <= simple_obj_ref_306_load_0_req_1;
      simple_obj_ref_379_load_0_ack_1 <= ackR(2);
      simple_obj_ref_282_load_0_ack_1 <= ackR(1);
      simple_obj_ref_306_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_379_word_address_0 & simple_obj_ref_282_word_address_0 & simple_obj_ref_306_word_address_0;
      simple_obj_ref_379_data_0 <= data_out(95 downto 64);
      simple_obj_ref_282_data_0 <= data_out(63 downto 32);
      simple_obj_ref_306_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 3,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(1),
          mack => memory_space_2_lr_ack(1),
          maddr => memory_space_2_lr_addr(1 downto 1),
          mtag => memory_space_2_lr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 3,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(1),
          mack => memory_space_2_lc_ack(1),
          mdata => memory_space_2_lc_data(63 downto 32),
          mtag => memory_space_2_lc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    -- shared load operator group (9) : simple_obj_ref_289_load_0 
    LoadGroup9: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_289_load_0_req_0;
      simple_obj_ref_289_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_289_load_0_req_1;
      simple_obj_ref_289_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_289_word_address_0;
      simple_obj_ref_289_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 9
    -- shared store operator group (0) : ptr_deref_223_store_0 ptr_deref_156_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_223_store_0_req_0;
      reqL(0) <= ptr_deref_156_store_0_req_0;
      ptr_deref_223_store_0_ack_0 <= ackL(1);
      ptr_deref_156_store_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_223_store_0_req_1;
      reqR(0) <= ptr_deref_156_store_0_req_1;
      ptr_deref_223_store_0_ack_1 <= ackR(1);
      ptr_deref_156_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_223_word_address_0 & ptr_deref_156_word_address_0;
      data_in <= ptr_deref_223_data_0 & ptr_deref_156_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_11_sr_req(0),
          mack => memory_space_11_sr_ack(0),
          maddr => memory_space_11_sr_addr(0 downto 0),
          mdata => memory_space_11_sr_data(31 downto 0),
          mtag => memory_space_11_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_11_sc_req(0),
          mack => memory_space_11_sc_ack(0),
          mtag => memory_space_11_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_210_store_0 ptr_deref_391_store_0 ptr_deref_235_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(8 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_210_store_0_req_0;
      reqL(1) <= ptr_deref_391_store_0_req_0;
      reqL(0) <= ptr_deref_235_store_0_req_0;
      ptr_deref_210_store_0_ack_0 <= ackL(2);
      ptr_deref_391_store_0_ack_0 <= ackL(1);
      ptr_deref_235_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_210_store_0_req_1;
      reqR(1) <= ptr_deref_391_store_0_req_1;
      reqR(0) <= ptr_deref_235_store_0_req_1;
      ptr_deref_210_store_0_ack_1 <= ackR(2);
      ptr_deref_391_store_0_ack_1 <= ackR(1);
      ptr_deref_235_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_210_word_address_0 & ptr_deref_391_word_address_0 & ptr_deref_235_word_address_0;
      data_in <= ptr_deref_210_data_0 & ptr_deref_391_data_0 & ptr_deref_235_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(2 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_258_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_258_store_0_req_0;
      ptr_deref_258_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_258_store_0_req_1;
      ptr_deref_258_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_258_word_address_0;
      data_in <= ptr_deref_258_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_12_sr_req(0),
          mack => memory_space_12_sr_ack(0),
          maddr => memory_space_12_sr_addr(0 downto 0),
          mdata => memory_space_12_sr_data(7 downto 0),
          mtag => memory_space_12_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_12_sc_req(0),
          mack => memory_space_12_sc_ack(0),
          mtag => memory_space_12_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_285_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_285_store_0_req_0;
      ptr_deref_285_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_285_store_0_req_1;
      ptr_deref_285_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_285_word_address_0;
      data_in <= ptr_deref_285_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_13_sr_req(0),
          mack => memory_space_13_sr_ack(0),
          maddr => memory_space_13_sr_addr(0 downto 0),
          mdata => memory_space_13_sr_data(31 downto 0),
          mtag => memory_space_13_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_13_sc_req(0),
          mack => memory_space_13_sc_ack(0),
          mtag => memory_space_13_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_375_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_375_store_0_req_0;
      ptr_deref_375_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_375_store_0_req_1;
      ptr_deref_375_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_375_word_address_0;
      data_in <= ptr_deref_375_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_14_sr_req(0),
          mack => memory_space_14_sr_ack(0),
          maddr => memory_space_14_sr_addr(0 downto 0),
          mdata => memory_space_14_sr_data(31 downto 0),
          mtag => memory_space_14_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_14_sc_req(0),
          mack => memory_space_14_sc_ack(0),
          mtag => memory_space_14_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : simple_obj_ref_317_store_0 simple_obj_ref_398_store_0 simple_obj_ref_243_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= simple_obj_ref_317_store_0_req_0;
      reqL(1) <= simple_obj_ref_398_store_0_req_0;
      reqL(0) <= simple_obj_ref_243_store_0_req_0;
      simple_obj_ref_317_store_0_ack_0 <= ackL(2);
      simple_obj_ref_398_store_0_ack_0 <= ackL(1);
      simple_obj_ref_243_store_0_ack_0 <= ackL(0);
      reqR(2) <= simple_obj_ref_317_store_0_req_1;
      reqR(1) <= simple_obj_ref_398_store_0_req_1;
      reqR(0) <= simple_obj_ref_243_store_0_req_1;
      simple_obj_ref_317_store_0_ack_1 <= ackR(2);
      simple_obj_ref_398_store_0_ack_1 <= ackR(1);
      simple_obj_ref_243_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_317_word_address_0 & simple_obj_ref_398_word_address_0 & simple_obj_ref_243_word_address_0;
      data_in <= simple_obj_ref_317_data_0 & simple_obj_ref_398_data_0 & simple_obj_ref_243_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared inport operator group (0) : simple_obj_ref_254_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_254_inst_req_0;
      simple_obj_ref_254_inst_ack_0 <= ack(0);
      simple_obj_ref_254_wire <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_request_pipe_read_req(0),
          oack => free_queue_request_pipe_read_ack(0),
          odata => free_queue_request_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_367_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_367_inst_req_0;
      simple_obj_ref_367_inst_ack_0 <= ack(0);
      simple_obj_ref_367_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_put_pipe_read_req(0),
          oack => free_queue_put_pipe_read_ack(0),
          odata => free_queue_put_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_335_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_335_inst_req_0;
      simple_obj_ref_335_inst_ack_0 <= ack(0);
      data_in <= type_cast_337_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_get_pipe_write_req(0),
          oack => free_queue_get_pipe_write_ack(0),
          odata => free_queue_get_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  RegisterBank_memory_space_11: register_bank -- 
    generic map(-- 
      num_loads => 3,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_11_lr_addr,
      lr_req_in => memory_space_11_lr_req,
      lr_ack_out => memory_space_11_lr_ack,
      lr_tag_in => memory_space_11_lr_tag,
      lc_req_in => memory_space_11_lc_req,
      lc_ack_out => memory_space_11_lc_ack,
      lc_data_out => memory_space_11_lc_data,
      lc_tag_out => memory_space_11_lc_tag,
      sr_addr_in => memory_space_11_sr_addr,
      sr_data_in => memory_space_11_sr_data,
      sr_req_in => memory_space_11_sr_req,
      sr_ack_out => memory_space_11_sr_ack,
      sr_tag_in => memory_space_11_sr_tag,
      sc_req_in=> memory_space_11_sc_req,
      sc_ack_out => memory_space_11_sc_ack,
      sc_tag_out => memory_space_11_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_12: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_12_lr_addr,
      lr_req_in => memory_space_12_lr_req,
      lr_ack_out => memory_space_12_lr_ack,
      lr_tag_in => memory_space_12_lr_tag,
      lc_req_in => memory_space_12_lc_req,
      lc_ack_out => memory_space_12_lc_ack,
      lc_data_out => memory_space_12_lc_data,
      lc_tag_out => memory_space_12_lc_tag,
      sr_addr_in => memory_space_12_sr_addr,
      sr_data_in => memory_space_12_sr_data,
      sr_req_in => memory_space_12_sr_req,
      sr_ack_out => memory_space_12_sr_ack,
      sr_tag_in => memory_space_12_sr_tag,
      sc_req_in=> memory_space_12_sc_req,
      sc_ack_out => memory_space_12_sc_ack,
      sc_tag_out => memory_space_12_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_13: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_13_lr_addr,
      lr_req_in => memory_space_13_lr_req,
      lr_ack_out => memory_space_13_lr_ack,
      lr_tag_in => memory_space_13_lr_tag,
      lc_req_in => memory_space_13_lc_req,
      lc_ack_out => memory_space_13_lc_ack,
      lc_data_out => memory_space_13_lc_data,
      lc_tag_out => memory_space_13_lc_tag,
      sr_addr_in => memory_space_13_sr_addr,
      sr_data_in => memory_space_13_sr_data,
      sr_req_in => memory_space_13_sr_req,
      sr_ack_out => memory_space_13_sr_ack,
      sr_tag_in => memory_space_13_sr_tag,
      sc_req_in=> memory_space_13_sc_req,
      sc_ack_out => memory_space_13_sc_ack,
      sc_tag_out => memory_space_13_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_14: register_bank -- 
    generic map(-- 
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_14_lr_addr,
      lr_req_in => memory_space_14_lr_req,
      lr_ack_out => memory_space_14_lr_ack,
      lr_tag_in => memory_space_14_lr_tag,
      lc_req_in => memory_space_14_lc_req,
      lc_ack_out => memory_space_14_lc_ack,
      lc_data_out => memory_space_14_lc_data,
      lc_tag_out => memory_space_14_lc_tag,
      sr_addr_in => memory_space_14_sr_addr,
      sr_data_in => memory_space_14_sr_data,
      sr_req_in => memory_space_14_sr_req,
      sr_ack_out => memory_space_14_sr_ack,
      sr_tag_in => memory_space_14_sr_tag,
      sc_req_in=> memory_space_14_sc_req,
      sc_ack_out => memory_space_14_sc_ack,
      sc_tag_out => memory_space_14_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity input_module is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(2 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_data_pipe_read_data : in   std_logic_vector(31 downto 0);
    foo_in_pipe_write_req : out  std_logic_vector(0 downto 0);
    foo_in_pipe_write_ack : in   std_logic_vector(0 downto 0);
    foo_in_pipe_write_data : out  std_logic_vector(31 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity input_module;
architecture Default of input_module is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_494_load_0_ack_0 : boolean;
  signal ptr_deref_489_gather_scatter_req_0 : boolean;
  signal ptr_deref_494_gather_scatter_ack_0 : boolean;
  signal ptr_deref_477_load_0_ack_1 : boolean;
  signal ptr_deref_477_load_0_req_1 : boolean;
  signal ptr_deref_481_gather_scatter_req_0 : boolean;
  signal ptr_deref_489_store_0_ack_0 : boolean;
  signal binary_453_inst_ack_1 : boolean;
  signal ptr_deref_446_load_0_req_1 : boolean;
  signal binary_453_inst_req_1 : boolean;
  signal type_cast_507_inst_req_0 : boolean;
  signal if_stmt_455_branch_ack_1 : boolean;
  signal ptr_deref_477_load_0_ack_0 : boolean;
  signal ptr_deref_446_gather_scatter_ack_0 : boolean;
  signal ptr_deref_494_load_0_req_1 : boolean;
  signal array_obj_ref_486_base_resize_ack_0 : boolean;
  signal array_obj_ref_486_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_423_inst_ack_0 : boolean;
  signal type_cast_498_inst_req_0 : boolean;
  signal array_obj_ref_486_base_resize_req_0 : boolean;
  signal if_stmt_455_branch_req_0 : boolean;
  signal ptr_deref_481_load_0_ack_1 : boolean;
  signal simple_obj_ref_433_inst_ack_0 : boolean;
  signal if_stmt_455_branch_ack_0 : boolean;
  signal type_cast_450_inst_req_0 : boolean;
  signal ptr_deref_472_store_0_ack_0 : boolean;
  signal ptr_deref_472_store_0_req_0 : boolean;
  signal ptr_deref_477_load_0_req_0 : boolean;
  signal type_cast_438_inst_ack_0 : boolean;
  signal array_obj_ref_486_root_address_inst_req_1 : boolean;
  signal ptr_deref_481_load_0_req_1 : boolean;
  signal type_cast_438_inst_req_0 : boolean;
  signal ptr_deref_472_gather_scatter_ack_0 : boolean;
  signal ptr_deref_477_gather_scatter_req_0 : boolean;
  signal ptr_deref_477_gather_scatter_ack_0 : boolean;
  signal ptr_deref_446_load_0_req_0 : boolean;
  signal ptr_deref_441_store_0_ack_0 : boolean;
  signal simple_obj_ref_505_inst_req_0 : boolean;
  signal array_obj_ref_486_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_486_root_address_inst_ack_1 : boolean;
  signal ptr_deref_489_store_0_ack_1 : boolean;
  signal ptr_deref_446_load_0_ack_1 : boolean;
  signal ptr_deref_446_gather_scatter_req_0 : boolean;
  signal ptr_deref_489_store_0_req_0 : boolean;
  signal ptr_deref_472_gather_scatter_req_0 : boolean;
  signal binary_453_inst_ack_0 : boolean;
  signal simple_obj_ref_423_inst_req_0 : boolean;
  signal type_cast_434_inst_ack_0 : boolean;
  signal ptr_deref_481_load_0_ack_0 : boolean;
  signal binary_453_inst_req_0 : boolean;
  signal ptr_deref_489_root_address_inst_ack_0 : boolean;
  signal type_cast_450_inst_ack_0 : boolean;
  signal ptr_deref_489_root_address_inst_req_0 : boolean;
  signal type_cast_434_inst_req_0 : boolean;
  signal ptr_deref_481_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_486_final_reg_req_0 : boolean;
  signal simple_obj_ref_505_inst_ack_0 : boolean;
  signal ptr_deref_446_load_0_ack_0 : boolean;
  signal array_obj_ref_486_final_reg_ack_0 : boolean;
  signal simple_obj_ref_433_inst_req_0 : boolean;
  signal ptr_deref_489_gather_scatter_ack_0 : boolean;
  signal ptr_deref_441_store_0_ack_1 : boolean;
  signal simple_obj_ref_468_inst_req_0 : boolean;
  signal ptr_deref_481_load_0_req_0 : boolean;
  signal ptr_deref_494_load_0_ack_1 : boolean;
  signal simple_obj_ref_468_inst_ack_0 : boolean;
  signal type_cast_498_inst_ack_0 : boolean;
  signal type_cast_507_inst_ack_0 : boolean;
  signal ptr_deref_489_addr_0_req_0 : boolean;
  signal ptr_deref_441_store_0_req_0 : boolean;
  signal ptr_deref_472_store_0_req_1 : boolean;
  signal type_cast_469_inst_req_0 : boolean;
  signal ptr_deref_472_store_0_ack_1 : boolean;
  signal ptr_deref_494_gather_scatter_req_0 : boolean;
  signal type_cast_469_inst_ack_0 : boolean;
  signal ptr_deref_494_load_0_req_0 : boolean;
  signal ptr_deref_489_addr_0_ack_0 : boolean;
  signal ptr_deref_441_gather_scatter_req_0 : boolean;
  signal ptr_deref_489_base_resize_req_0 : boolean;
  signal ptr_deref_441_gather_scatter_ack_0 : boolean;
  signal ptr_deref_489_base_resize_ack_0 : boolean;
  signal ptr_deref_441_store_0_req_1 : boolean;
  signal ptr_deref_489_store_0_req_1 : boolean;
  signal memory_space_15_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_15_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_15_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_15_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_15_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_15_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_15_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_15_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_15_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_15_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_15_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_15_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_15_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_15_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_15_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_15_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_16_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_16_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_16_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_16_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_16_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_16_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_16_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_16_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_16_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_16_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_16_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_16_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_16_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_16_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_16_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_16_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  input_module_CP_1810: Block -- control-path 
    signal input_module_CP_1810_start: Boolean;
    signal Xentry_1811_symbol: Boolean;
    signal Xexit_1812_symbol: Boolean;
    signal branch_block_stmt_405_1813_symbol : Boolean;
    -- 
  begin -- 
    input_module_CP_1810_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_1811_symbol  <= input_module_CP_1810_start; -- transition $entry
    branch_block_stmt_405_1813: Block -- branch_block_stmt_405 
      signal branch_block_stmt_405_1813_start: Boolean;
      signal Xentry_1814_symbol: Boolean;
      signal Xexit_1815_symbol: Boolean;
      signal branch_block_stmt_405_x_xentry_x_xx_x1816_symbol : Boolean;
      signal branch_block_stmt_405_x_xexit_x_xx_x1817_symbol : Boolean;
      signal assign_stmt_411_to_assign_stmt_415_x_xentry_x_xx_x1818_symbol : Boolean;
      signal assign_stmt_411_to_assign_stmt_415_x_xexit_x_xx_x1819_symbol : Boolean;
      signal bb_0_bb_1_1820_symbol : Boolean;
      signal merge_stmt_417_x_xexit_x_xx_x1821_symbol : Boolean;
      signal assign_stmt_422_x_xentry_x_xx_x1822_symbol : Boolean;
      signal assign_stmt_422_x_xexit_x_xx_x1823_symbol : Boolean;
      signal assign_stmt_426_x_xentry_x_xx_x1824_symbol : Boolean;
      signal assign_stmt_426_x_xexit_x_xx_x1825_symbol : Boolean;
      signal assign_stmt_431_x_xentry_x_xx_x1826_symbol : Boolean;
      signal assign_stmt_431_x_xexit_x_xx_x1827_symbol : Boolean;
      signal assign_stmt_435_x_xentry_x_xx_x1828_symbol : Boolean;
      signal assign_stmt_435_x_xexit_x_xx_x1829_symbol : Boolean;
      signal assign_stmt_439_to_assign_stmt_454_x_xentry_x_xx_x1830_symbol : Boolean;
      signal assign_stmt_439_to_assign_stmt_454_x_xexit_x_xx_x1831_symbol : Boolean;
      signal if_stmt_455_x_xentry_x_xx_x1832_symbol : Boolean;
      signal if_stmt_455_x_xexit_x_xx_x1833_symbol : Boolean;
      signal merge_stmt_461_x_xentry_x_xx_x1834_symbol : Boolean;
      signal merge_stmt_461_x_xexit_x_xx_x1835_symbol : Boolean;
      signal assign_stmt_466_x_xentry_x_xx_x1836_symbol : Boolean;
      signal assign_stmt_466_x_xexit_x_xx_x1837_symbol : Boolean;
      signal assign_stmt_470_x_xentry_x_xx_x1838_symbol : Boolean;
      signal assign_stmt_470_x_xexit_x_xx_x1839_symbol : Boolean;
      signal assign_stmt_474_to_assign_stmt_504_x_xentry_x_xx_x1840_symbol : Boolean;
      signal assign_stmt_474_to_assign_stmt_504_x_xexit_x_xx_x1841_symbol : Boolean;
      signal assign_stmt_508_x_xentry_x_xx_x1842_symbol : Boolean;
      signal assign_stmt_508_x_xexit_x_xx_x1843_symbol : Boolean;
      signal bb_2_bb_1_1844_symbol : Boolean;
      signal assign_stmt_411_to_assign_stmt_415_1845_symbol : Boolean;
      signal assign_stmt_422_1848_symbol : Boolean;
      signal assign_stmt_426_1851_symbol : Boolean;
      signal assign_stmt_431_1862_symbol : Boolean;
      signal assign_stmt_435_1865_symbol : Boolean;
      signal assign_stmt_439_to_assign_stmt_454_1883_symbol : Boolean;
      signal if_stmt_455_dead_link_1978_symbol : Boolean;
      signal if_stmt_455_eval_test_1982_symbol : Boolean;
      signal simple_obj_ref_456_place_1986_symbol : Boolean;
      signal if_stmt_455_if_link_1987_symbol : Boolean;
      signal if_stmt_455_else_link_1991_symbol : Boolean;
      signal bb_1_bb_2_1995_symbol : Boolean;
      signal bb_1_bb_1_1996_symbol : Boolean;
      signal assign_stmt_466_1997_symbol : Boolean;
      signal assign_stmt_470_2000_symbol : Boolean;
      signal assign_stmt_474_to_assign_stmt_504_2018_symbol : Boolean;
      signal assign_stmt_508_2230_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_2249_symbol : Boolean;
      signal bb_1_bb_1_PhiReq_2252_symbol : Boolean;
      signal bb_2_bb_1_PhiReq_2255_symbol : Boolean;
      signal merge_stmt_417_PhiReqMerge_2258_symbol : Boolean;
      signal merge_stmt_417_PhiAck_2259_symbol : Boolean;
      signal merge_stmt_461_dead_link_2263_symbol : Boolean;
      signal bb_1_bb_2_PhiReq_2267_symbol : Boolean;
      signal merge_stmt_461_PhiReqMerge_2270_symbol : Boolean;
      signal merge_stmt_461_PhiAck_2271_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_405_1813_start <= Xentry_1811_symbol; -- control passed to block
      Xentry_1814_symbol  <= branch_block_stmt_405_1813_start; -- transition branch_block_stmt_405/$entry
      branch_block_stmt_405_x_xentry_x_xx_x1816_symbol  <=  Xentry_1814_symbol; -- place branch_block_stmt_405/branch_block_stmt_405__entry__ (optimized away) 
      branch_block_stmt_405_x_xexit_x_xx_x1817_symbol  <=   false ; -- place branch_block_stmt_405/branch_block_stmt_405__exit__ (optimized away) 
      assign_stmt_411_to_assign_stmt_415_x_xentry_x_xx_x1818_symbol  <=  branch_block_stmt_405_x_xentry_x_xx_x1816_symbol; -- place branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415__entry__ (optimized away) 
      assign_stmt_411_to_assign_stmt_415_x_xexit_x_xx_x1819_symbol  <=  assign_stmt_411_to_assign_stmt_415_1845_symbol; -- place branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415__exit__ (optimized away) 
      bb_0_bb_1_1820_symbol  <=  assign_stmt_411_to_assign_stmt_415_x_xexit_x_xx_x1819_symbol; -- place branch_block_stmt_405/bb_0_bb_1 (optimized away) 
      merge_stmt_417_x_xexit_x_xx_x1821_symbol  <=  merge_stmt_417_PhiAck_2259_symbol; -- place branch_block_stmt_405/merge_stmt_417__exit__ (optimized away) 
      assign_stmt_422_x_xentry_x_xx_x1822_symbol  <=  merge_stmt_417_x_xexit_x_xx_x1821_symbol; -- place branch_block_stmt_405/assign_stmt_422__entry__ (optimized away) 
      assign_stmt_422_x_xexit_x_xx_x1823_symbol  <=  assign_stmt_422_1848_symbol; -- place branch_block_stmt_405/assign_stmt_422__exit__ (optimized away) 
      assign_stmt_426_x_xentry_x_xx_x1824_symbol  <=  assign_stmt_422_x_xexit_x_xx_x1823_symbol; -- place branch_block_stmt_405/assign_stmt_426__entry__ (optimized away) 
      assign_stmt_426_x_xexit_x_xx_x1825_symbol  <=  assign_stmt_426_1851_symbol; -- place branch_block_stmt_405/assign_stmt_426__exit__ (optimized away) 
      assign_stmt_431_x_xentry_x_xx_x1826_symbol  <=  assign_stmt_426_x_xexit_x_xx_x1825_symbol; -- place branch_block_stmt_405/assign_stmt_431__entry__ (optimized away) 
      assign_stmt_431_x_xexit_x_xx_x1827_symbol  <=  assign_stmt_431_1862_symbol; -- place branch_block_stmt_405/assign_stmt_431__exit__ (optimized away) 
      assign_stmt_435_x_xentry_x_xx_x1828_symbol  <=  assign_stmt_431_x_xexit_x_xx_x1827_symbol; -- place branch_block_stmt_405/assign_stmt_435__entry__ (optimized away) 
      assign_stmt_435_x_xexit_x_xx_x1829_symbol  <=  assign_stmt_435_1865_symbol; -- place branch_block_stmt_405/assign_stmt_435__exit__ (optimized away) 
      assign_stmt_439_to_assign_stmt_454_x_xentry_x_xx_x1830_symbol  <=  assign_stmt_435_x_xexit_x_xx_x1829_symbol; -- place branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454__entry__ (optimized away) 
      assign_stmt_439_to_assign_stmt_454_x_xexit_x_xx_x1831_symbol  <=  assign_stmt_439_to_assign_stmt_454_1883_symbol; -- place branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454__exit__ (optimized away) 
      if_stmt_455_x_xentry_x_xx_x1832_symbol  <=  assign_stmt_439_to_assign_stmt_454_x_xexit_x_xx_x1831_symbol; -- place branch_block_stmt_405/if_stmt_455__entry__ (optimized away) 
      if_stmt_455_x_xexit_x_xx_x1833_symbol  <=  if_stmt_455_dead_link_1978_symbol; -- place branch_block_stmt_405/if_stmt_455__exit__ (optimized away) 
      merge_stmt_461_x_xentry_x_xx_x1834_symbol  <=  if_stmt_455_x_xexit_x_xx_x1833_symbol; -- place branch_block_stmt_405/merge_stmt_461__entry__ (optimized away) 
      merge_stmt_461_x_xexit_x_xx_x1835_symbol  <=  merge_stmt_461_dead_link_2263_symbol or merge_stmt_461_PhiAck_2271_symbol; -- place branch_block_stmt_405/merge_stmt_461__exit__ (optimized away) 
      assign_stmt_466_x_xentry_x_xx_x1836_symbol  <=  merge_stmt_461_x_xexit_x_xx_x1835_symbol; -- place branch_block_stmt_405/assign_stmt_466__entry__ (optimized away) 
      assign_stmt_466_x_xexit_x_xx_x1837_symbol  <=  assign_stmt_466_1997_symbol; -- place branch_block_stmt_405/assign_stmt_466__exit__ (optimized away) 
      assign_stmt_470_x_xentry_x_xx_x1838_symbol  <=  assign_stmt_466_x_xexit_x_xx_x1837_symbol; -- place branch_block_stmt_405/assign_stmt_470__entry__ (optimized away) 
      assign_stmt_470_x_xexit_x_xx_x1839_symbol  <=  assign_stmt_470_2000_symbol; -- place branch_block_stmt_405/assign_stmt_470__exit__ (optimized away) 
      assign_stmt_474_to_assign_stmt_504_x_xentry_x_xx_x1840_symbol  <=  assign_stmt_470_x_xexit_x_xx_x1839_symbol; -- place branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504__entry__ (optimized away) 
      assign_stmt_474_to_assign_stmt_504_x_xexit_x_xx_x1841_symbol  <=  assign_stmt_474_to_assign_stmt_504_2018_symbol; -- place branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504__exit__ (optimized away) 
      assign_stmt_508_x_xentry_x_xx_x1842_symbol  <=  assign_stmt_474_to_assign_stmt_504_x_xexit_x_xx_x1841_symbol; -- place branch_block_stmt_405/assign_stmt_508__entry__ (optimized away) 
      assign_stmt_508_x_xexit_x_xx_x1843_symbol  <=  assign_stmt_508_2230_symbol; -- place branch_block_stmt_405/assign_stmt_508__exit__ (optimized away) 
      bb_2_bb_1_1844_symbol  <=  assign_stmt_508_x_xexit_x_xx_x1843_symbol; -- place branch_block_stmt_405/bb_2_bb_1 (optimized away) 
      assign_stmt_411_to_assign_stmt_415_1845: Block -- branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415 
        signal assign_stmt_411_to_assign_stmt_415_1845_start: Boolean;
        signal Xentry_1846_symbol: Boolean;
        signal Xexit_1847_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_411_to_assign_stmt_415_1845_start <= assign_stmt_411_to_assign_stmt_415_x_xentry_x_xx_x1818_symbol; -- control passed to block
        Xentry_1846_symbol  <= assign_stmt_411_to_assign_stmt_415_1845_start; -- transition branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415/$entry
        Xexit_1847_symbol <= Xentry_1846_symbol; -- transition branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415/$exit
        assign_stmt_411_to_assign_stmt_415_1845_symbol <= Xexit_1847_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_411_to_assign_stmt_415
      assign_stmt_422_1848: Block -- branch_block_stmt_405/assign_stmt_422 
        signal assign_stmt_422_1848_start: Boolean;
        signal Xentry_1849_symbol: Boolean;
        signal Xexit_1850_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_422_1848_start <= assign_stmt_422_x_xentry_x_xx_x1822_symbol; -- control passed to block
        Xentry_1849_symbol  <= assign_stmt_422_1848_start; -- transition branch_block_stmt_405/assign_stmt_422/$entry
        Xexit_1850_symbol <= Xentry_1849_symbol; -- transition branch_block_stmt_405/assign_stmt_422/$exit
        assign_stmt_422_1848_symbol <= Xexit_1850_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_422
      assign_stmt_426_1851: Block -- branch_block_stmt_405/assign_stmt_426 
        signal assign_stmt_426_1851_start: Boolean;
        signal Xentry_1852_symbol: Boolean;
        signal Xexit_1853_symbol: Boolean;
        signal assign_stmt_426_active_x_x1854_symbol : Boolean;
        signal assign_stmt_426_completed_x_x1855_symbol : Boolean;
        signal simple_obj_ref_423_trigger_x_x1856_symbol : Boolean;
        signal simple_obj_ref_423_complete_1857_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_426_1851_start <= assign_stmt_426_x_xentry_x_xx_x1824_symbol; -- control passed to block
        Xentry_1852_symbol  <= assign_stmt_426_1851_start; -- transition branch_block_stmt_405/assign_stmt_426/$entry
        assign_stmt_426_active_x_x1854_symbol <= Xentry_1852_symbol; -- transition branch_block_stmt_405/assign_stmt_426/assign_stmt_426_active_
        assign_stmt_426_completed_x_x1855_symbol <= simple_obj_ref_423_complete_1857_symbol; -- transition branch_block_stmt_405/assign_stmt_426/assign_stmt_426_completed_
        simple_obj_ref_423_trigger_x_x1856_symbol <= assign_stmt_426_active_x_x1854_symbol; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_trigger_
        simple_obj_ref_423_complete_1857: Block -- branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete 
          signal simple_obj_ref_423_complete_1857_start: Boolean;
          signal Xentry_1858_symbol: Boolean;
          signal Xexit_1859_symbol: Boolean;
          signal pipe_wreq_1860_symbol : Boolean;
          signal pipe_wack_1861_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_423_complete_1857_start <= simple_obj_ref_423_trigger_x_x1856_symbol; -- control passed to block
          Xentry_1858_symbol  <= simple_obj_ref_423_complete_1857_start; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/$entry
          pipe_wreq_1860_symbol <= Xentry_1858_symbol; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/pipe_wreq
          simple_obj_ref_423_inst_req_0 <= pipe_wreq_1860_symbol; -- link to DP
          pipe_wack_1861_symbol <= simple_obj_ref_423_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/pipe_wack
          Xexit_1859_symbol <= pipe_wack_1861_symbol; -- transition branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete/$exit
          simple_obj_ref_423_complete_1857_symbol <= Xexit_1859_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_426/simple_obj_ref_423_complete
        Xexit_1853_symbol <= assign_stmt_426_completed_x_x1855_symbol; -- transition branch_block_stmt_405/assign_stmt_426/$exit
        assign_stmt_426_1851_symbol <= Xexit_1853_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_426
      assign_stmt_431_1862: Block -- branch_block_stmt_405/assign_stmt_431 
        signal assign_stmt_431_1862_start: Boolean;
        signal Xentry_1863_symbol: Boolean;
        signal Xexit_1864_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_431_1862_start <= assign_stmt_431_x_xentry_x_xx_x1826_symbol; -- control passed to block
        Xentry_1863_symbol  <= assign_stmt_431_1862_start; -- transition branch_block_stmt_405/assign_stmt_431/$entry
        Xexit_1864_symbol <= Xentry_1863_symbol; -- transition branch_block_stmt_405/assign_stmt_431/$exit
        assign_stmt_431_1862_symbol <= Xexit_1864_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_431
      assign_stmt_435_1865: Block -- branch_block_stmt_405/assign_stmt_435 
        signal assign_stmt_435_1865_start: Boolean;
        signal Xentry_1866_symbol: Boolean;
        signal Xexit_1867_symbol: Boolean;
        signal assign_stmt_435_active_x_x1868_symbol : Boolean;
        signal assign_stmt_435_completed_x_x1869_symbol : Boolean;
        signal type_cast_434_active_x_x1870_symbol : Boolean;
        signal type_cast_434_trigger_x_x1871_symbol : Boolean;
        signal simple_obj_ref_433_trigger_x_x1872_symbol : Boolean;
        signal simple_obj_ref_433_complete_1873_symbol : Boolean;
        signal type_cast_434_complete_1878_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_435_1865_start <= assign_stmt_435_x_xentry_x_xx_x1828_symbol; -- control passed to block
        Xentry_1866_symbol  <= assign_stmt_435_1865_start; -- transition branch_block_stmt_405/assign_stmt_435/$entry
        assign_stmt_435_active_x_x1868_symbol <= type_cast_434_complete_1878_symbol; -- transition branch_block_stmt_405/assign_stmt_435/assign_stmt_435_active_
        assign_stmt_435_completed_x_x1869_symbol <= assign_stmt_435_active_x_x1868_symbol; -- transition branch_block_stmt_405/assign_stmt_435/assign_stmt_435_completed_
        type_cast_434_active_x_x1870_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_435/type_cast_434_active_ 
          signal type_cast_434_active_x_x1870_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_434_active_x_x1870_predecessors(0) <= type_cast_434_trigger_x_x1871_symbol;
          type_cast_434_active_x_x1870_predecessors(1) <= simple_obj_ref_433_complete_1873_symbol;
          type_cast_434_active_x_x1870_join: join -- 
            port map( -- 
              preds => type_cast_434_active_x_x1870_predecessors,
              symbol_out => type_cast_434_active_x_x1870_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_435/type_cast_434_active_
        type_cast_434_trigger_x_x1871_symbol <= Xentry_1866_symbol; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_trigger_
        simple_obj_ref_433_trigger_x_x1872_symbol <= Xentry_1866_symbol; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_trigger_
        simple_obj_ref_433_complete_1873: Block -- branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete 
          signal simple_obj_ref_433_complete_1873_start: Boolean;
          signal Xentry_1874_symbol: Boolean;
          signal Xexit_1875_symbol: Boolean;
          signal req_1876_symbol : Boolean;
          signal ack_1877_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_433_complete_1873_start <= simple_obj_ref_433_trigger_x_x1872_symbol; -- control passed to block
          Xentry_1874_symbol  <= simple_obj_ref_433_complete_1873_start; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/$entry
          req_1876_symbol <= Xentry_1874_symbol; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/req
          simple_obj_ref_433_inst_req_0 <= req_1876_symbol; -- link to DP
          ack_1877_symbol <= simple_obj_ref_433_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/ack
          Xexit_1875_symbol <= ack_1877_symbol; -- transition branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete/$exit
          simple_obj_ref_433_complete_1873_symbol <= Xexit_1875_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_435/simple_obj_ref_433_complete
        type_cast_434_complete_1878: Block -- branch_block_stmt_405/assign_stmt_435/type_cast_434_complete 
          signal type_cast_434_complete_1878_start: Boolean;
          signal Xentry_1879_symbol: Boolean;
          signal Xexit_1880_symbol: Boolean;
          signal req_1881_symbol : Boolean;
          signal ack_1882_symbol : Boolean;
          -- 
        begin -- 
          type_cast_434_complete_1878_start <= type_cast_434_active_x_x1870_symbol; -- control passed to block
          Xentry_1879_symbol  <= type_cast_434_complete_1878_start; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/$entry
          req_1881_symbol <= Xentry_1879_symbol; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/req
          type_cast_434_inst_req_0 <= req_1881_symbol; -- link to DP
          ack_1882_symbol <= type_cast_434_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/ack
          Xexit_1880_symbol <= ack_1882_symbol; -- transition branch_block_stmt_405/assign_stmt_435/type_cast_434_complete/$exit
          type_cast_434_complete_1878_symbol <= Xexit_1880_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_435/type_cast_434_complete
        Xexit_1867_symbol <= assign_stmt_435_completed_x_x1869_symbol; -- transition branch_block_stmt_405/assign_stmt_435/$exit
        assign_stmt_435_1865_symbol <= Xexit_1867_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_435
      assign_stmt_439_to_assign_stmt_454_1883: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454 
        signal assign_stmt_439_to_assign_stmt_454_1883_start: Boolean;
        signal Xentry_1884_symbol: Boolean;
        signal Xexit_1885_symbol: Boolean;
        signal assign_stmt_439_active_x_x1886_symbol : Boolean;
        signal assign_stmt_439_completed_x_x1887_symbol : Boolean;
        signal type_cast_438_active_x_x1888_symbol : Boolean;
        signal type_cast_438_trigger_x_x1889_symbol : Boolean;
        signal simple_obj_ref_437_complete_1890_symbol : Boolean;
        signal type_cast_438_complete_1891_symbol : Boolean;
        signal assign_stmt_443_active_x_x1896_symbol : Boolean;
        signal assign_stmt_443_completed_x_x1897_symbol : Boolean;
        signal simple_obj_ref_442_complete_1898_symbol : Boolean;
        signal ptr_deref_441_trigger_x_x1899_symbol : Boolean;
        signal ptr_deref_441_active_x_x1900_symbol : Boolean;
        signal ptr_deref_441_base_address_calculated_1901_symbol : Boolean;
        signal ptr_deref_441_root_address_calculated_1902_symbol : Boolean;
        signal ptr_deref_441_word_address_calculated_1903_symbol : Boolean;
        signal ptr_deref_441_request_1904_symbol : Boolean;
        signal ptr_deref_441_complete_1917_symbol : Boolean;
        signal assign_stmt_447_active_x_x1928_symbol : Boolean;
        signal assign_stmt_447_completed_x_x1929_symbol : Boolean;
        signal ptr_deref_446_trigger_x_x1930_symbol : Boolean;
        signal ptr_deref_446_active_x_x1931_symbol : Boolean;
        signal ptr_deref_446_base_address_calculated_1932_symbol : Boolean;
        signal ptr_deref_446_root_address_calculated_1933_symbol : Boolean;
        signal ptr_deref_446_word_address_calculated_1934_symbol : Boolean;
        signal ptr_deref_446_request_1935_symbol : Boolean;
        signal ptr_deref_446_complete_1946_symbol : Boolean;
        signal assign_stmt_454_active_x_x1959_symbol : Boolean;
        signal assign_stmt_454_completed_x_x1960_symbol : Boolean;
        signal binary_453_active_x_x1961_symbol : Boolean;
        signal binary_453_trigger_x_x1962_symbol : Boolean;
        signal type_cast_450_active_x_x1963_symbol : Boolean;
        signal type_cast_450_trigger_x_x1964_symbol : Boolean;
        signal simple_obj_ref_449_complete_1965_symbol : Boolean;
        signal type_cast_450_complete_1966_symbol : Boolean;
        signal binary_453_complete_1971_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_439_to_assign_stmt_454_1883_start <= assign_stmt_439_to_assign_stmt_454_x_xentry_x_xx_x1830_symbol; -- control passed to block
        Xentry_1884_symbol  <= assign_stmt_439_to_assign_stmt_454_1883_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/$entry
        assign_stmt_439_active_x_x1886_symbol <= type_cast_438_complete_1891_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_439_active_
        assign_stmt_439_completed_x_x1887_symbol <= assign_stmt_439_active_x_x1886_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_439_completed_
        type_cast_438_active_x_x1888_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_active_ 
          signal type_cast_438_active_x_x1888_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_438_active_x_x1888_predecessors(0) <= type_cast_438_trigger_x_x1889_symbol;
          type_cast_438_active_x_x1888_predecessors(1) <= simple_obj_ref_437_complete_1890_symbol;
          type_cast_438_active_x_x1888_join: join -- 
            port map( -- 
              preds => type_cast_438_active_x_x1888_predecessors,
              symbol_out => type_cast_438_active_x_x1888_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_active_
        type_cast_438_trigger_x_x1889_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_trigger_
        simple_obj_ref_437_complete_1890_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/simple_obj_ref_437_complete
        type_cast_438_complete_1891: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete 
          signal type_cast_438_complete_1891_start: Boolean;
          signal Xentry_1892_symbol: Boolean;
          signal Xexit_1893_symbol: Boolean;
          signal req_1894_symbol : Boolean;
          signal ack_1895_symbol : Boolean;
          -- 
        begin -- 
          type_cast_438_complete_1891_start <= type_cast_438_active_x_x1888_symbol; -- control passed to block
          Xentry_1892_symbol  <= type_cast_438_complete_1891_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/$entry
          req_1894_symbol <= Xentry_1892_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/req
          type_cast_438_inst_req_0 <= req_1894_symbol; -- link to DP
          ack_1895_symbol <= type_cast_438_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/ack
          Xexit_1893_symbol <= ack_1895_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete/$exit
          type_cast_438_complete_1891_symbol <= Xexit_1893_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_438_complete
        assign_stmt_443_active_x_x1896_symbol <= simple_obj_ref_442_complete_1898_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_443_active_
        assign_stmt_443_completed_x_x1897_symbol <= ptr_deref_441_complete_1917_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_443_completed_
        simple_obj_ref_442_complete_1898_symbol <= assign_stmt_439_completed_x_x1887_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/simple_obj_ref_442_complete
        ptr_deref_441_trigger_x_x1899_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_trigger_ 
          signal ptr_deref_441_trigger_x_x1899_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_441_trigger_x_x1899_predecessors(0) <= ptr_deref_441_word_address_calculated_1903_symbol;
          ptr_deref_441_trigger_x_x1899_predecessors(1) <= assign_stmt_443_active_x_x1896_symbol;
          ptr_deref_441_trigger_x_x1899_join: join -- 
            port map( -- 
              preds => ptr_deref_441_trigger_x_x1899_predecessors,
              symbol_out => ptr_deref_441_trigger_x_x1899_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_trigger_
        ptr_deref_441_active_x_x1900_symbol <= ptr_deref_441_request_1904_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_active_
        ptr_deref_441_base_address_calculated_1901_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_base_address_calculated
        ptr_deref_441_root_address_calculated_1902_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_root_address_calculated
        ptr_deref_441_word_address_calculated_1903_symbol <= ptr_deref_441_root_address_calculated_1902_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_word_address_calculated
        ptr_deref_441_request_1904: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request 
          signal ptr_deref_441_request_1904_start: Boolean;
          signal Xentry_1905_symbol: Boolean;
          signal Xexit_1906_symbol: Boolean;
          signal split_req_1907_symbol : Boolean;
          signal split_ack_1908_symbol : Boolean;
          signal word_access_1909_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_441_request_1904_start <= ptr_deref_441_trigger_x_x1899_symbol; -- control passed to block
          Xentry_1905_symbol  <= ptr_deref_441_request_1904_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/$entry
          split_req_1907_symbol <= Xentry_1905_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/split_req
          ptr_deref_441_gather_scatter_req_0 <= split_req_1907_symbol; -- link to DP
          split_ack_1908_symbol <= ptr_deref_441_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/split_ack
          word_access_1909: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access 
            signal word_access_1909_start: Boolean;
            signal Xentry_1910_symbol: Boolean;
            signal Xexit_1911_symbol: Boolean;
            signal word_access_0_1912_symbol : Boolean;
            -- 
          begin -- 
            word_access_1909_start <= split_ack_1908_symbol; -- control passed to block
            Xentry_1910_symbol  <= word_access_1909_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/$entry
            word_access_0_1912: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0 
              signal word_access_0_1912_start: Boolean;
              signal Xentry_1913_symbol: Boolean;
              signal Xexit_1914_symbol: Boolean;
              signal rr_1915_symbol : Boolean;
              signal ra_1916_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1912_start <= Xentry_1910_symbol; -- control passed to block
              Xentry_1913_symbol  <= word_access_0_1912_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/$entry
              rr_1915_symbol <= Xentry_1913_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/rr
              ptr_deref_441_store_0_req_0 <= rr_1915_symbol; -- link to DP
              ra_1916_symbol <= ptr_deref_441_store_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/ra
              Xexit_1914_symbol <= ra_1916_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0/$exit
              word_access_0_1912_symbol <= Xexit_1914_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/word_access_0
            Xexit_1911_symbol <= word_access_0_1912_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access/$exit
            word_access_1909_symbol <= Xexit_1911_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/word_access
          Xexit_1906_symbol <= word_access_1909_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request/$exit
          ptr_deref_441_request_1904_symbol <= Xexit_1906_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_request
        ptr_deref_441_complete_1917: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete 
          signal ptr_deref_441_complete_1917_start: Boolean;
          signal Xentry_1918_symbol: Boolean;
          signal Xexit_1919_symbol: Boolean;
          signal word_access_1920_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_441_complete_1917_start <= ptr_deref_441_active_x_x1900_symbol; -- control passed to block
          Xentry_1918_symbol  <= ptr_deref_441_complete_1917_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/$entry
          word_access_1920: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access 
            signal word_access_1920_start: Boolean;
            signal Xentry_1921_symbol: Boolean;
            signal Xexit_1922_symbol: Boolean;
            signal word_access_0_1923_symbol : Boolean;
            -- 
          begin -- 
            word_access_1920_start <= Xentry_1918_symbol; -- control passed to block
            Xentry_1921_symbol  <= word_access_1920_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/$entry
            word_access_0_1923: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0 
              signal word_access_0_1923_start: Boolean;
              signal Xentry_1924_symbol: Boolean;
              signal Xexit_1925_symbol: Boolean;
              signal cr_1926_symbol : Boolean;
              signal ca_1927_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1923_start <= Xentry_1921_symbol; -- control passed to block
              Xentry_1924_symbol  <= word_access_0_1923_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/$entry
              cr_1926_symbol <= Xentry_1924_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/cr
              ptr_deref_441_store_0_req_1 <= cr_1926_symbol; -- link to DP
              ca_1927_symbol <= ptr_deref_441_store_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/ca
              Xexit_1925_symbol <= ca_1927_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0/$exit
              word_access_0_1923_symbol <= Xexit_1925_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/word_access_0
            Xexit_1922_symbol <= word_access_0_1923_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access/$exit
            word_access_1920_symbol <= Xexit_1922_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/word_access
          Xexit_1919_symbol <= word_access_1920_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete/$exit
          ptr_deref_441_complete_1917_symbol <= Xexit_1919_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_441_complete
        assign_stmt_447_active_x_x1928_symbol <= ptr_deref_446_complete_1946_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_447_active_
        assign_stmt_447_completed_x_x1929_symbol <= assign_stmt_447_active_x_x1928_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_447_completed_
        ptr_deref_446_trigger_x_x1930_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_trigger_ 
          signal ptr_deref_446_trigger_x_x1930_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_446_trigger_x_x1930_predecessors(0) <= ptr_deref_446_word_address_calculated_1934_symbol;
          ptr_deref_446_trigger_x_x1930_predecessors(1) <= ptr_deref_441_active_x_x1900_symbol;
          ptr_deref_446_trigger_x_x1930_join: join -- 
            port map( -- 
              preds => ptr_deref_446_trigger_x_x1930_predecessors,
              symbol_out => ptr_deref_446_trigger_x_x1930_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_trigger_
        ptr_deref_446_active_x_x1931_symbol <= ptr_deref_446_request_1935_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_active_
        ptr_deref_446_base_address_calculated_1932_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_base_address_calculated
        ptr_deref_446_root_address_calculated_1933_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_root_address_calculated
        ptr_deref_446_word_address_calculated_1934_symbol <= ptr_deref_446_root_address_calculated_1933_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_word_address_calculated
        ptr_deref_446_request_1935: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request 
          signal ptr_deref_446_request_1935_start: Boolean;
          signal Xentry_1936_symbol: Boolean;
          signal Xexit_1937_symbol: Boolean;
          signal word_access_1938_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_446_request_1935_start <= ptr_deref_446_trigger_x_x1930_symbol; -- control passed to block
          Xentry_1936_symbol  <= ptr_deref_446_request_1935_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/$entry
          word_access_1938: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access 
            signal word_access_1938_start: Boolean;
            signal Xentry_1939_symbol: Boolean;
            signal Xexit_1940_symbol: Boolean;
            signal word_access_0_1941_symbol : Boolean;
            -- 
          begin -- 
            word_access_1938_start <= Xentry_1936_symbol; -- control passed to block
            Xentry_1939_symbol  <= word_access_1938_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/$entry
            word_access_0_1941: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0 
              signal word_access_0_1941_start: Boolean;
              signal Xentry_1942_symbol: Boolean;
              signal Xexit_1943_symbol: Boolean;
              signal rr_1944_symbol : Boolean;
              signal ra_1945_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1941_start <= Xentry_1939_symbol; -- control passed to block
              Xentry_1942_symbol  <= word_access_0_1941_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/$entry
              rr_1944_symbol <= Xentry_1942_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/rr
              ptr_deref_446_load_0_req_0 <= rr_1944_symbol; -- link to DP
              ra_1945_symbol <= ptr_deref_446_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/ra
              Xexit_1943_symbol <= ra_1945_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0/$exit
              word_access_0_1941_symbol <= Xexit_1943_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/word_access_0
            Xexit_1940_symbol <= word_access_0_1941_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access/$exit
            word_access_1938_symbol <= Xexit_1940_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/word_access
          Xexit_1937_symbol <= word_access_1938_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request/$exit
          ptr_deref_446_request_1935_symbol <= Xexit_1937_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_request
        ptr_deref_446_complete_1946: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete 
          signal ptr_deref_446_complete_1946_start: Boolean;
          signal Xentry_1947_symbol: Boolean;
          signal Xexit_1948_symbol: Boolean;
          signal word_access_1949_symbol : Boolean;
          signal merge_req_1957_symbol : Boolean;
          signal merge_ack_1958_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_446_complete_1946_start <= ptr_deref_446_active_x_x1931_symbol; -- control passed to block
          Xentry_1947_symbol  <= ptr_deref_446_complete_1946_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/$entry
          word_access_1949: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access 
            signal word_access_1949_start: Boolean;
            signal Xentry_1950_symbol: Boolean;
            signal Xexit_1951_symbol: Boolean;
            signal word_access_0_1952_symbol : Boolean;
            -- 
          begin -- 
            word_access_1949_start <= Xentry_1947_symbol; -- control passed to block
            Xentry_1950_symbol  <= word_access_1949_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/$entry
            word_access_0_1952: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0 
              signal word_access_0_1952_start: Boolean;
              signal Xentry_1953_symbol: Boolean;
              signal Xexit_1954_symbol: Boolean;
              signal cr_1955_symbol : Boolean;
              signal ca_1956_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_1952_start <= Xentry_1950_symbol; -- control passed to block
              Xentry_1953_symbol  <= word_access_0_1952_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/$entry
              cr_1955_symbol <= Xentry_1953_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/cr
              ptr_deref_446_load_0_req_1 <= cr_1955_symbol; -- link to DP
              ca_1956_symbol <= ptr_deref_446_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/ca
              Xexit_1954_symbol <= ca_1956_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0/$exit
              word_access_0_1952_symbol <= Xexit_1954_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/word_access_0
            Xexit_1951_symbol <= word_access_0_1952_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access/$exit
            word_access_1949_symbol <= Xexit_1951_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/word_access
          merge_req_1957_symbol <= word_access_1949_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/merge_req
          ptr_deref_446_gather_scatter_req_0 <= merge_req_1957_symbol; -- link to DP
          merge_ack_1958_symbol <= ptr_deref_446_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/merge_ack
          Xexit_1948_symbol <= merge_ack_1958_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete/$exit
          ptr_deref_446_complete_1946_symbol <= Xexit_1948_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/ptr_deref_446_complete
        assign_stmt_454_active_x_x1959_symbol <= binary_453_complete_1971_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_454_active_
        assign_stmt_454_completed_x_x1960_symbol <= assign_stmt_454_active_x_x1959_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/assign_stmt_454_completed_
        binary_453_active_x_x1961_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_active_ 
          signal binary_453_active_x_x1961_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          binary_453_active_x_x1961_predecessors(0) <= binary_453_trigger_x_x1962_symbol;
          binary_453_active_x_x1961_predecessors(1) <= type_cast_450_complete_1966_symbol;
          binary_453_active_x_x1961_join: join -- 
            port map( -- 
              preds => binary_453_active_x_x1961_predecessors,
              symbol_out => binary_453_active_x_x1961_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_active_
        binary_453_trigger_x_x1962_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_trigger_
        type_cast_450_active_x_x1963_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_active_ 
          signal type_cast_450_active_x_x1963_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_450_active_x_x1963_predecessors(0) <= type_cast_450_trigger_x_x1964_symbol;
          type_cast_450_active_x_x1963_predecessors(1) <= simple_obj_ref_449_complete_1965_symbol;
          type_cast_450_active_x_x1963_join: join -- 
            port map( -- 
              preds => type_cast_450_active_x_x1963_predecessors,
              symbol_out => type_cast_450_active_x_x1963_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_active_
        type_cast_450_trigger_x_x1964_symbol <= Xentry_1884_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_trigger_
        simple_obj_ref_449_complete_1965_symbol <= assign_stmt_447_completed_x_x1929_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/simple_obj_ref_449_complete
        type_cast_450_complete_1966: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete 
          signal type_cast_450_complete_1966_start: Boolean;
          signal Xentry_1967_symbol: Boolean;
          signal Xexit_1968_symbol: Boolean;
          signal req_1969_symbol : Boolean;
          signal ack_1970_symbol : Boolean;
          -- 
        begin -- 
          type_cast_450_complete_1966_start <= type_cast_450_active_x_x1963_symbol; -- control passed to block
          Xentry_1967_symbol  <= type_cast_450_complete_1966_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/$entry
          req_1969_symbol <= Xentry_1967_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/req
          type_cast_450_inst_req_0 <= req_1969_symbol; -- link to DP
          ack_1970_symbol <= type_cast_450_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/ack
          Xexit_1968_symbol <= ack_1970_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete/$exit
          type_cast_450_complete_1966_symbol <= Xexit_1968_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/type_cast_450_complete
        binary_453_complete_1971: Block -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete 
          signal binary_453_complete_1971_start: Boolean;
          signal Xentry_1972_symbol: Boolean;
          signal Xexit_1973_symbol: Boolean;
          signal rr_1974_symbol : Boolean;
          signal ra_1975_symbol : Boolean;
          signal cr_1976_symbol : Boolean;
          signal ca_1977_symbol : Boolean;
          -- 
        begin -- 
          binary_453_complete_1971_start <= binary_453_active_x_x1961_symbol; -- control passed to block
          Xentry_1972_symbol  <= binary_453_complete_1971_start; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/$entry
          rr_1974_symbol <= Xentry_1972_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/rr
          binary_453_inst_req_0 <= rr_1974_symbol; -- link to DP
          ra_1975_symbol <= binary_453_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/ra
          cr_1976_symbol <= ra_1975_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/cr
          binary_453_inst_req_1 <= cr_1976_symbol; -- link to DP
          ca_1977_symbol <= binary_453_inst_ack_1; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/ca
          Xexit_1973_symbol <= ca_1977_symbol; -- transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete/$exit
          binary_453_complete_1971_symbol <= Xexit_1973_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/binary_453_complete
        Xexit_1885_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/$exit 
          signal Xexit_1885_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          Xexit_1885_predecessors(0) <= assign_stmt_443_completed_x_x1897_symbol;
          Xexit_1885_predecessors(1) <= ptr_deref_441_base_address_calculated_1901_symbol;
          Xexit_1885_predecessors(2) <= ptr_deref_446_base_address_calculated_1932_symbol;
          Xexit_1885_predecessors(3) <= assign_stmt_454_completed_x_x1960_symbol;
          Xexit_1885_join: join -- 
            port map( -- 
              preds => Xexit_1885_predecessors,
              symbol_out => Xexit_1885_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454/$exit
        assign_stmt_439_to_assign_stmt_454_1883_symbol <= Xexit_1885_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_439_to_assign_stmt_454
      if_stmt_455_dead_link_1978: Block -- branch_block_stmt_405/if_stmt_455_dead_link 
        signal if_stmt_455_dead_link_1978_start: Boolean;
        signal Xentry_1979_symbol: Boolean;
        signal Xexit_1980_symbol: Boolean;
        signal dead_transition_1981_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_dead_link_1978_start <= if_stmt_455_x_xentry_x_xx_x1832_symbol; -- control passed to block
        Xentry_1979_symbol  <= if_stmt_455_dead_link_1978_start; -- transition branch_block_stmt_405/if_stmt_455_dead_link/$entry
        dead_transition_1981_symbol <= false;
        Xexit_1980_symbol <= dead_transition_1981_symbol; -- transition branch_block_stmt_405/if_stmt_455_dead_link/$exit
        if_stmt_455_dead_link_1978_symbol <= Xexit_1980_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_dead_link
      if_stmt_455_eval_test_1982: Block -- branch_block_stmt_405/if_stmt_455_eval_test 
        signal if_stmt_455_eval_test_1982_start: Boolean;
        signal Xentry_1983_symbol: Boolean;
        signal Xexit_1984_symbol: Boolean;
        signal branch_req_1985_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_eval_test_1982_start <= if_stmt_455_x_xentry_x_xx_x1832_symbol; -- control passed to block
        Xentry_1983_symbol  <= if_stmt_455_eval_test_1982_start; -- transition branch_block_stmt_405/if_stmt_455_eval_test/$entry
        branch_req_1985_symbol <= Xentry_1983_symbol; -- transition branch_block_stmt_405/if_stmt_455_eval_test/branch_req
        if_stmt_455_branch_req_0 <= branch_req_1985_symbol; -- link to DP
        Xexit_1984_symbol <= branch_req_1985_symbol; -- transition branch_block_stmt_405/if_stmt_455_eval_test/$exit
        if_stmt_455_eval_test_1982_symbol <= Xexit_1984_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_eval_test
      simple_obj_ref_456_place_1986_symbol  <=  if_stmt_455_eval_test_1982_symbol; -- place branch_block_stmt_405/simple_obj_ref_456_place (optimized away) 
      if_stmt_455_if_link_1987: Block -- branch_block_stmt_405/if_stmt_455_if_link 
        signal if_stmt_455_if_link_1987_start: Boolean;
        signal Xentry_1988_symbol: Boolean;
        signal Xexit_1989_symbol: Boolean;
        signal if_choice_transition_1990_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_if_link_1987_start <= simple_obj_ref_456_place_1986_symbol; -- control passed to block
        Xentry_1988_symbol  <= if_stmt_455_if_link_1987_start; -- transition branch_block_stmt_405/if_stmt_455_if_link/$entry
        if_choice_transition_1990_symbol <= if_stmt_455_branch_ack_1; -- transition branch_block_stmt_405/if_stmt_455_if_link/if_choice_transition
        Xexit_1989_symbol <= if_choice_transition_1990_symbol; -- transition branch_block_stmt_405/if_stmt_455_if_link/$exit
        if_stmt_455_if_link_1987_symbol <= Xexit_1989_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_if_link
      if_stmt_455_else_link_1991: Block -- branch_block_stmt_405/if_stmt_455_else_link 
        signal if_stmt_455_else_link_1991_start: Boolean;
        signal Xentry_1992_symbol: Boolean;
        signal Xexit_1993_symbol: Boolean;
        signal else_choice_transition_1994_symbol : Boolean;
        -- 
      begin -- 
        if_stmt_455_else_link_1991_start <= simple_obj_ref_456_place_1986_symbol; -- control passed to block
        Xentry_1992_symbol  <= if_stmt_455_else_link_1991_start; -- transition branch_block_stmt_405/if_stmt_455_else_link/$entry
        else_choice_transition_1994_symbol <= if_stmt_455_branch_ack_0; -- transition branch_block_stmt_405/if_stmt_455_else_link/else_choice_transition
        Xexit_1993_symbol <= else_choice_transition_1994_symbol; -- transition branch_block_stmt_405/if_stmt_455_else_link/$exit
        if_stmt_455_else_link_1991_symbol <= Xexit_1993_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/if_stmt_455_else_link
      bb_1_bb_2_1995_symbol  <=  if_stmt_455_if_link_1987_symbol; -- place branch_block_stmt_405/bb_1_bb_2 (optimized away) 
      bb_1_bb_1_1996_symbol  <=  if_stmt_455_else_link_1991_symbol; -- place branch_block_stmt_405/bb_1_bb_1 (optimized away) 
      assign_stmt_466_1997: Block -- branch_block_stmt_405/assign_stmt_466 
        signal assign_stmt_466_1997_start: Boolean;
        signal Xentry_1998_symbol: Boolean;
        signal Xexit_1999_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_466_1997_start <= assign_stmt_466_x_xentry_x_xx_x1836_symbol; -- control passed to block
        Xentry_1998_symbol  <= assign_stmt_466_1997_start; -- transition branch_block_stmt_405/assign_stmt_466/$entry
        Xexit_1999_symbol <= Xentry_1998_symbol; -- transition branch_block_stmt_405/assign_stmt_466/$exit
        assign_stmt_466_1997_symbol <= Xexit_1999_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_466
      assign_stmt_470_2000: Block -- branch_block_stmt_405/assign_stmt_470 
        signal assign_stmt_470_2000_start: Boolean;
        signal Xentry_2001_symbol: Boolean;
        signal Xexit_2002_symbol: Boolean;
        signal assign_stmt_470_active_x_x2003_symbol : Boolean;
        signal assign_stmt_470_completed_x_x2004_symbol : Boolean;
        signal type_cast_469_active_x_x2005_symbol : Boolean;
        signal type_cast_469_trigger_x_x2006_symbol : Boolean;
        signal simple_obj_ref_468_trigger_x_x2007_symbol : Boolean;
        signal simple_obj_ref_468_complete_2008_symbol : Boolean;
        signal type_cast_469_complete_2013_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_470_2000_start <= assign_stmt_470_x_xentry_x_xx_x1838_symbol; -- control passed to block
        Xentry_2001_symbol  <= assign_stmt_470_2000_start; -- transition branch_block_stmt_405/assign_stmt_470/$entry
        assign_stmt_470_active_x_x2003_symbol <= type_cast_469_complete_2013_symbol; -- transition branch_block_stmt_405/assign_stmt_470/assign_stmt_470_active_
        assign_stmt_470_completed_x_x2004_symbol <= assign_stmt_470_active_x_x2003_symbol; -- transition branch_block_stmt_405/assign_stmt_470/assign_stmt_470_completed_
        type_cast_469_active_x_x2005_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_470/type_cast_469_active_ 
          signal type_cast_469_active_x_x2005_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_469_active_x_x2005_predecessors(0) <= type_cast_469_trigger_x_x2006_symbol;
          type_cast_469_active_x_x2005_predecessors(1) <= simple_obj_ref_468_complete_2008_symbol;
          type_cast_469_active_x_x2005_join: join -- 
            port map( -- 
              preds => type_cast_469_active_x_x2005_predecessors,
              symbol_out => type_cast_469_active_x_x2005_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_470/type_cast_469_active_
        type_cast_469_trigger_x_x2006_symbol <= Xentry_2001_symbol; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_trigger_
        simple_obj_ref_468_trigger_x_x2007_symbol <= Xentry_2001_symbol; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_trigger_
        simple_obj_ref_468_complete_2008: Block -- branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete 
          signal simple_obj_ref_468_complete_2008_start: Boolean;
          signal Xentry_2009_symbol: Boolean;
          signal Xexit_2010_symbol: Boolean;
          signal req_2011_symbol : Boolean;
          signal ack_2012_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_468_complete_2008_start <= simple_obj_ref_468_trigger_x_x2007_symbol; -- control passed to block
          Xentry_2009_symbol  <= simple_obj_ref_468_complete_2008_start; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/$entry
          req_2011_symbol <= Xentry_2009_symbol; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/req
          simple_obj_ref_468_inst_req_0 <= req_2011_symbol; -- link to DP
          ack_2012_symbol <= simple_obj_ref_468_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/ack
          Xexit_2010_symbol <= ack_2012_symbol; -- transition branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete/$exit
          simple_obj_ref_468_complete_2008_symbol <= Xexit_2010_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_470/simple_obj_ref_468_complete
        type_cast_469_complete_2013: Block -- branch_block_stmt_405/assign_stmt_470/type_cast_469_complete 
          signal type_cast_469_complete_2013_start: Boolean;
          signal Xentry_2014_symbol: Boolean;
          signal Xexit_2015_symbol: Boolean;
          signal req_2016_symbol : Boolean;
          signal ack_2017_symbol : Boolean;
          -- 
        begin -- 
          type_cast_469_complete_2013_start <= type_cast_469_active_x_x2005_symbol; -- control passed to block
          Xentry_2014_symbol  <= type_cast_469_complete_2013_start; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/$entry
          req_2016_symbol <= Xentry_2014_symbol; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/req
          type_cast_469_inst_req_0 <= req_2016_symbol; -- link to DP
          ack_2017_symbol <= type_cast_469_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/ack
          Xexit_2015_symbol <= ack_2017_symbol; -- transition branch_block_stmt_405/assign_stmt_470/type_cast_469_complete/$exit
          type_cast_469_complete_2013_symbol <= Xexit_2015_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_470/type_cast_469_complete
        Xexit_2002_symbol <= assign_stmt_470_completed_x_x2004_symbol; -- transition branch_block_stmt_405/assign_stmt_470/$exit
        assign_stmt_470_2000_symbol <= Xexit_2002_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_470
      assign_stmt_474_to_assign_stmt_504_2018: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504 
        signal assign_stmt_474_to_assign_stmt_504_2018_start: Boolean;
        signal Xentry_2019_symbol: Boolean;
        signal Xexit_2020_symbol: Boolean;
        signal assign_stmt_474_active_x_x2021_symbol : Boolean;
        signal assign_stmt_474_completed_x_x2022_symbol : Boolean;
        signal simple_obj_ref_473_complete_2023_symbol : Boolean;
        signal ptr_deref_472_trigger_x_x2024_symbol : Boolean;
        signal ptr_deref_472_active_x_x2025_symbol : Boolean;
        signal ptr_deref_472_base_address_calculated_2026_symbol : Boolean;
        signal ptr_deref_472_root_address_calculated_2027_symbol : Boolean;
        signal ptr_deref_472_word_address_calculated_2028_symbol : Boolean;
        signal ptr_deref_472_request_2029_symbol : Boolean;
        signal ptr_deref_472_complete_2042_symbol : Boolean;
        signal assign_stmt_478_active_x_x2053_symbol : Boolean;
        signal assign_stmt_478_completed_x_x2054_symbol : Boolean;
        signal ptr_deref_477_trigger_x_x2055_symbol : Boolean;
        signal ptr_deref_477_active_x_x2056_symbol : Boolean;
        signal ptr_deref_477_base_address_calculated_2057_symbol : Boolean;
        signal ptr_deref_477_root_address_calculated_2058_symbol : Boolean;
        signal ptr_deref_477_word_address_calculated_2059_symbol : Boolean;
        signal ptr_deref_477_request_2060_symbol : Boolean;
        signal ptr_deref_477_complete_2071_symbol : Boolean;
        signal assign_stmt_482_active_x_x2084_symbol : Boolean;
        signal assign_stmt_482_completed_x_x2085_symbol : Boolean;
        signal ptr_deref_481_trigger_x_x2086_symbol : Boolean;
        signal ptr_deref_481_active_x_x2087_symbol : Boolean;
        signal ptr_deref_481_base_address_calculated_2088_symbol : Boolean;
        signal ptr_deref_481_root_address_calculated_2089_symbol : Boolean;
        signal ptr_deref_481_word_address_calculated_2090_symbol : Boolean;
        signal ptr_deref_481_request_2091_symbol : Boolean;
        signal ptr_deref_481_complete_2102_symbol : Boolean;
        signal assign_stmt_487_active_x_x2115_symbol : Boolean;
        signal assign_stmt_487_completed_x_x2116_symbol : Boolean;
        signal array_obj_ref_486_trigger_x_x2117_symbol : Boolean;
        signal array_obj_ref_486_active_x_x2118_symbol : Boolean;
        signal array_obj_ref_486_base_address_calculated_2119_symbol : Boolean;
        signal array_obj_ref_486_root_address_calculated_2120_symbol : Boolean;
        signal array_obj_ref_486_base_address_resized_2121_symbol : Boolean;
        signal array_obj_ref_486_base_addr_resize_2122_symbol : Boolean;
        signal array_obj_ref_486_base_plus_offset_trigger_2127_symbol : Boolean;
        signal array_obj_ref_486_base_plus_offset_2128_symbol : Boolean;
        signal array_obj_ref_486_complete_2135_symbol : Boolean;
        signal assign_stmt_491_active_x_x2140_symbol : Boolean;
        signal assign_stmt_491_completed_x_x2141_symbol : Boolean;
        signal simple_obj_ref_490_complete_2142_symbol : Boolean;
        signal ptr_deref_489_trigger_x_x2143_symbol : Boolean;
        signal ptr_deref_489_active_x_x2144_symbol : Boolean;
        signal ptr_deref_489_base_address_calculated_2145_symbol : Boolean;
        signal simple_obj_ref_488_complete_2146_symbol : Boolean;
        signal ptr_deref_489_root_address_calculated_2147_symbol : Boolean;
        signal ptr_deref_489_word_address_calculated_2148_symbol : Boolean;
        signal ptr_deref_489_base_address_resized_2149_symbol : Boolean;
        signal ptr_deref_489_base_addr_resize_2150_symbol : Boolean;
        signal ptr_deref_489_base_plus_offset_2155_symbol : Boolean;
        signal ptr_deref_489_word_addrgen_2160_symbol : Boolean;
        signal ptr_deref_489_request_2165_symbol : Boolean;
        signal ptr_deref_489_complete_2178_symbol : Boolean;
        signal assign_stmt_495_active_x_x2189_symbol : Boolean;
        signal assign_stmt_495_completed_x_x2190_symbol : Boolean;
        signal ptr_deref_494_trigger_x_x2191_symbol : Boolean;
        signal ptr_deref_494_active_x_x2192_symbol : Boolean;
        signal ptr_deref_494_base_address_calculated_2193_symbol : Boolean;
        signal ptr_deref_494_root_address_calculated_2194_symbol : Boolean;
        signal ptr_deref_494_word_address_calculated_2195_symbol : Boolean;
        signal ptr_deref_494_request_2196_symbol : Boolean;
        signal ptr_deref_494_complete_2207_symbol : Boolean;
        signal assign_stmt_499_active_x_x2220_symbol : Boolean;
        signal assign_stmt_499_completed_x_x2221_symbol : Boolean;
        signal type_cast_498_active_x_x2222_symbol : Boolean;
        signal type_cast_498_trigger_x_x2223_symbol : Boolean;
        signal simple_obj_ref_497_complete_2224_symbol : Boolean;
        signal type_cast_498_complete_2225_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_474_to_assign_stmt_504_2018_start <= assign_stmt_474_to_assign_stmt_504_x_xentry_x_xx_x1840_symbol; -- control passed to block
        Xentry_2019_symbol  <= assign_stmt_474_to_assign_stmt_504_2018_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/$entry
        assign_stmt_474_active_x_x2021_symbol <= simple_obj_ref_473_complete_2023_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_474_active_
        assign_stmt_474_completed_x_x2022_symbol <= ptr_deref_472_complete_2042_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_474_completed_
        simple_obj_ref_473_complete_2023_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_473_complete
        ptr_deref_472_trigger_x_x2024_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_trigger_ 
          signal ptr_deref_472_trigger_x_x2024_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_472_trigger_x_x2024_predecessors(0) <= ptr_deref_472_word_address_calculated_2028_symbol;
          ptr_deref_472_trigger_x_x2024_predecessors(1) <= assign_stmt_474_active_x_x2021_symbol;
          ptr_deref_472_trigger_x_x2024_join: join -- 
            port map( -- 
              preds => ptr_deref_472_trigger_x_x2024_predecessors,
              symbol_out => ptr_deref_472_trigger_x_x2024_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_trigger_
        ptr_deref_472_active_x_x2025_symbol <= ptr_deref_472_request_2029_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_active_
        ptr_deref_472_base_address_calculated_2026_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_base_address_calculated
        ptr_deref_472_root_address_calculated_2027_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_root_address_calculated
        ptr_deref_472_word_address_calculated_2028_symbol <= ptr_deref_472_root_address_calculated_2027_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_word_address_calculated
        ptr_deref_472_request_2029: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request 
          signal ptr_deref_472_request_2029_start: Boolean;
          signal Xentry_2030_symbol: Boolean;
          signal Xexit_2031_symbol: Boolean;
          signal split_req_2032_symbol : Boolean;
          signal split_ack_2033_symbol : Boolean;
          signal word_access_2034_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_472_request_2029_start <= ptr_deref_472_trigger_x_x2024_symbol; -- control passed to block
          Xentry_2030_symbol  <= ptr_deref_472_request_2029_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/$entry
          split_req_2032_symbol <= Xentry_2030_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/split_req
          ptr_deref_472_gather_scatter_req_0 <= split_req_2032_symbol; -- link to DP
          split_ack_2033_symbol <= ptr_deref_472_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/split_ack
          word_access_2034: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access 
            signal word_access_2034_start: Boolean;
            signal Xentry_2035_symbol: Boolean;
            signal Xexit_2036_symbol: Boolean;
            signal word_access_0_2037_symbol : Boolean;
            -- 
          begin -- 
            word_access_2034_start <= split_ack_2033_symbol; -- control passed to block
            Xentry_2035_symbol  <= word_access_2034_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/$entry
            word_access_0_2037: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0 
              signal word_access_0_2037_start: Boolean;
              signal Xentry_2038_symbol: Boolean;
              signal Xexit_2039_symbol: Boolean;
              signal rr_2040_symbol : Boolean;
              signal ra_2041_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2037_start <= Xentry_2035_symbol; -- control passed to block
              Xentry_2038_symbol  <= word_access_0_2037_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/$entry
              rr_2040_symbol <= Xentry_2038_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/rr
              ptr_deref_472_store_0_req_0 <= rr_2040_symbol; -- link to DP
              ra_2041_symbol <= ptr_deref_472_store_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/ra
              Xexit_2039_symbol <= ra_2041_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0/$exit
              word_access_0_2037_symbol <= Xexit_2039_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/word_access_0
            Xexit_2036_symbol <= word_access_0_2037_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access/$exit
            word_access_2034_symbol <= Xexit_2036_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/word_access
          Xexit_2031_symbol <= word_access_2034_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request/$exit
          ptr_deref_472_request_2029_symbol <= Xexit_2031_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_request
        ptr_deref_472_complete_2042: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete 
          signal ptr_deref_472_complete_2042_start: Boolean;
          signal Xentry_2043_symbol: Boolean;
          signal Xexit_2044_symbol: Boolean;
          signal word_access_2045_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_472_complete_2042_start <= ptr_deref_472_active_x_x2025_symbol; -- control passed to block
          Xentry_2043_symbol  <= ptr_deref_472_complete_2042_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/$entry
          word_access_2045: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access 
            signal word_access_2045_start: Boolean;
            signal Xentry_2046_symbol: Boolean;
            signal Xexit_2047_symbol: Boolean;
            signal word_access_0_2048_symbol : Boolean;
            -- 
          begin -- 
            word_access_2045_start <= Xentry_2043_symbol; -- control passed to block
            Xentry_2046_symbol  <= word_access_2045_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/$entry
            word_access_0_2048: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0 
              signal word_access_0_2048_start: Boolean;
              signal Xentry_2049_symbol: Boolean;
              signal Xexit_2050_symbol: Boolean;
              signal cr_2051_symbol : Boolean;
              signal ca_2052_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2048_start <= Xentry_2046_symbol; -- control passed to block
              Xentry_2049_symbol  <= word_access_0_2048_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/$entry
              cr_2051_symbol <= Xentry_2049_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/cr
              ptr_deref_472_store_0_req_1 <= cr_2051_symbol; -- link to DP
              ca_2052_symbol <= ptr_deref_472_store_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/ca
              Xexit_2050_symbol <= ca_2052_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0/$exit
              word_access_0_2048_symbol <= Xexit_2050_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/word_access_0
            Xexit_2047_symbol <= word_access_0_2048_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access/$exit
            word_access_2045_symbol <= Xexit_2047_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/word_access
          Xexit_2044_symbol <= word_access_2045_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete/$exit
          ptr_deref_472_complete_2042_symbol <= Xexit_2044_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_472_complete
        assign_stmt_478_active_x_x2053_symbol <= ptr_deref_477_complete_2071_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_478_active_
        assign_stmt_478_completed_x_x2054_symbol <= assign_stmt_478_active_x_x2053_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_478_completed_
        ptr_deref_477_trigger_x_x2055_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_trigger_ 
          signal ptr_deref_477_trigger_x_x2055_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_477_trigger_x_x2055_predecessors(0) <= ptr_deref_477_word_address_calculated_2059_symbol;
          ptr_deref_477_trigger_x_x2055_predecessors(1) <= ptr_deref_472_active_x_x2025_symbol;
          ptr_deref_477_trigger_x_x2055_join: join -- 
            port map( -- 
              preds => ptr_deref_477_trigger_x_x2055_predecessors,
              symbol_out => ptr_deref_477_trigger_x_x2055_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_trigger_
        ptr_deref_477_active_x_x2056_symbol <= ptr_deref_477_request_2060_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_active_
        ptr_deref_477_base_address_calculated_2057_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_base_address_calculated
        ptr_deref_477_root_address_calculated_2058_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_root_address_calculated
        ptr_deref_477_word_address_calculated_2059_symbol <= ptr_deref_477_root_address_calculated_2058_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_word_address_calculated
        ptr_deref_477_request_2060: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request 
          signal ptr_deref_477_request_2060_start: Boolean;
          signal Xentry_2061_symbol: Boolean;
          signal Xexit_2062_symbol: Boolean;
          signal word_access_2063_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_477_request_2060_start <= ptr_deref_477_trigger_x_x2055_symbol; -- control passed to block
          Xentry_2061_symbol  <= ptr_deref_477_request_2060_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/$entry
          word_access_2063: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access 
            signal word_access_2063_start: Boolean;
            signal Xentry_2064_symbol: Boolean;
            signal Xexit_2065_symbol: Boolean;
            signal word_access_0_2066_symbol : Boolean;
            -- 
          begin -- 
            word_access_2063_start <= Xentry_2061_symbol; -- control passed to block
            Xentry_2064_symbol  <= word_access_2063_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/$entry
            word_access_0_2066: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0 
              signal word_access_0_2066_start: Boolean;
              signal Xentry_2067_symbol: Boolean;
              signal Xexit_2068_symbol: Boolean;
              signal rr_2069_symbol : Boolean;
              signal ra_2070_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2066_start <= Xentry_2064_symbol; -- control passed to block
              Xentry_2067_symbol  <= word_access_0_2066_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/$entry
              rr_2069_symbol <= Xentry_2067_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/rr
              ptr_deref_477_load_0_req_0 <= rr_2069_symbol; -- link to DP
              ra_2070_symbol <= ptr_deref_477_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/ra
              Xexit_2068_symbol <= ra_2070_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0/$exit
              word_access_0_2066_symbol <= Xexit_2068_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/word_access_0
            Xexit_2065_symbol <= word_access_0_2066_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access/$exit
            word_access_2063_symbol <= Xexit_2065_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/word_access
          Xexit_2062_symbol <= word_access_2063_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request/$exit
          ptr_deref_477_request_2060_symbol <= Xexit_2062_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_request
        ptr_deref_477_complete_2071: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete 
          signal ptr_deref_477_complete_2071_start: Boolean;
          signal Xentry_2072_symbol: Boolean;
          signal Xexit_2073_symbol: Boolean;
          signal word_access_2074_symbol : Boolean;
          signal merge_req_2082_symbol : Boolean;
          signal merge_ack_2083_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_477_complete_2071_start <= ptr_deref_477_active_x_x2056_symbol; -- control passed to block
          Xentry_2072_symbol  <= ptr_deref_477_complete_2071_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/$entry
          word_access_2074: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access 
            signal word_access_2074_start: Boolean;
            signal Xentry_2075_symbol: Boolean;
            signal Xexit_2076_symbol: Boolean;
            signal word_access_0_2077_symbol : Boolean;
            -- 
          begin -- 
            word_access_2074_start <= Xentry_2072_symbol; -- control passed to block
            Xentry_2075_symbol  <= word_access_2074_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/$entry
            word_access_0_2077: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0 
              signal word_access_0_2077_start: Boolean;
              signal Xentry_2078_symbol: Boolean;
              signal Xexit_2079_symbol: Boolean;
              signal cr_2080_symbol : Boolean;
              signal ca_2081_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2077_start <= Xentry_2075_symbol; -- control passed to block
              Xentry_2078_symbol  <= word_access_0_2077_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/$entry
              cr_2080_symbol <= Xentry_2078_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/cr
              ptr_deref_477_load_0_req_1 <= cr_2080_symbol; -- link to DP
              ca_2081_symbol <= ptr_deref_477_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/ca
              Xexit_2079_symbol <= ca_2081_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0/$exit
              word_access_0_2077_symbol <= Xexit_2079_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/word_access_0
            Xexit_2076_symbol <= word_access_0_2077_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access/$exit
            word_access_2074_symbol <= Xexit_2076_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/word_access
          merge_req_2082_symbol <= word_access_2074_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/merge_req
          ptr_deref_477_gather_scatter_req_0 <= merge_req_2082_symbol; -- link to DP
          merge_ack_2083_symbol <= ptr_deref_477_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/merge_ack
          Xexit_2073_symbol <= merge_ack_2083_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete/$exit
          ptr_deref_477_complete_2071_symbol <= Xexit_2073_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_477_complete
        assign_stmt_482_active_x_x2084_symbol <= ptr_deref_481_complete_2102_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_482_active_
        assign_stmt_482_completed_x_x2085_symbol <= assign_stmt_482_active_x_x2084_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_482_completed_
        ptr_deref_481_trigger_x_x2086_symbol <= ptr_deref_481_word_address_calculated_2090_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_trigger_
        ptr_deref_481_active_x_x2087_symbol <= ptr_deref_481_request_2091_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_active_
        ptr_deref_481_base_address_calculated_2088_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_base_address_calculated
        ptr_deref_481_root_address_calculated_2089_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_root_address_calculated
        ptr_deref_481_word_address_calculated_2090_symbol <= ptr_deref_481_root_address_calculated_2089_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_word_address_calculated
        ptr_deref_481_request_2091: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request 
          signal ptr_deref_481_request_2091_start: Boolean;
          signal Xentry_2092_symbol: Boolean;
          signal Xexit_2093_symbol: Boolean;
          signal word_access_2094_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_481_request_2091_start <= ptr_deref_481_trigger_x_x2086_symbol; -- control passed to block
          Xentry_2092_symbol  <= ptr_deref_481_request_2091_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/$entry
          word_access_2094: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access 
            signal word_access_2094_start: Boolean;
            signal Xentry_2095_symbol: Boolean;
            signal Xexit_2096_symbol: Boolean;
            signal word_access_0_2097_symbol : Boolean;
            -- 
          begin -- 
            word_access_2094_start <= Xentry_2092_symbol; -- control passed to block
            Xentry_2095_symbol  <= word_access_2094_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/$entry
            word_access_0_2097: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0 
              signal word_access_0_2097_start: Boolean;
              signal Xentry_2098_symbol: Boolean;
              signal Xexit_2099_symbol: Boolean;
              signal rr_2100_symbol : Boolean;
              signal ra_2101_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2097_start <= Xentry_2095_symbol; -- control passed to block
              Xentry_2098_symbol  <= word_access_0_2097_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/$entry
              rr_2100_symbol <= Xentry_2098_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/rr
              ptr_deref_481_load_0_req_0 <= rr_2100_symbol; -- link to DP
              ra_2101_symbol <= ptr_deref_481_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/ra
              Xexit_2099_symbol <= ra_2101_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0/$exit
              word_access_0_2097_symbol <= Xexit_2099_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/word_access_0
            Xexit_2096_symbol <= word_access_0_2097_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access/$exit
            word_access_2094_symbol <= Xexit_2096_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/word_access
          Xexit_2093_symbol <= word_access_2094_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request/$exit
          ptr_deref_481_request_2091_symbol <= Xexit_2093_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_request
        ptr_deref_481_complete_2102: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete 
          signal ptr_deref_481_complete_2102_start: Boolean;
          signal Xentry_2103_symbol: Boolean;
          signal Xexit_2104_symbol: Boolean;
          signal word_access_2105_symbol : Boolean;
          signal merge_req_2113_symbol : Boolean;
          signal merge_ack_2114_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_481_complete_2102_start <= ptr_deref_481_active_x_x2087_symbol; -- control passed to block
          Xentry_2103_symbol  <= ptr_deref_481_complete_2102_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/$entry
          word_access_2105: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access 
            signal word_access_2105_start: Boolean;
            signal Xentry_2106_symbol: Boolean;
            signal Xexit_2107_symbol: Boolean;
            signal word_access_0_2108_symbol : Boolean;
            -- 
          begin -- 
            word_access_2105_start <= Xentry_2103_symbol; -- control passed to block
            Xentry_2106_symbol  <= word_access_2105_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/$entry
            word_access_0_2108: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0 
              signal word_access_0_2108_start: Boolean;
              signal Xentry_2109_symbol: Boolean;
              signal Xexit_2110_symbol: Boolean;
              signal cr_2111_symbol : Boolean;
              signal ca_2112_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2108_start <= Xentry_2106_symbol; -- control passed to block
              Xentry_2109_symbol  <= word_access_0_2108_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/$entry
              cr_2111_symbol <= Xentry_2109_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/cr
              ptr_deref_481_load_0_req_1 <= cr_2111_symbol; -- link to DP
              ca_2112_symbol <= ptr_deref_481_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/ca
              Xexit_2110_symbol <= ca_2112_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0/$exit
              word_access_0_2108_symbol <= Xexit_2110_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/word_access_0
            Xexit_2107_symbol <= word_access_0_2108_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access/$exit
            word_access_2105_symbol <= Xexit_2107_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/word_access
          merge_req_2113_symbol <= word_access_2105_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/merge_req
          ptr_deref_481_gather_scatter_req_0 <= merge_req_2113_symbol; -- link to DP
          merge_ack_2114_symbol <= ptr_deref_481_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/merge_ack
          Xexit_2104_symbol <= merge_ack_2114_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete/$exit
          ptr_deref_481_complete_2102_symbol <= Xexit_2104_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_481_complete
        assign_stmt_487_active_x_x2115_symbol <= array_obj_ref_486_complete_2135_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_487_active_
        assign_stmt_487_completed_x_x2116_symbol <= assign_stmt_487_active_x_x2115_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_487_completed_
        array_obj_ref_486_trigger_x_x2117_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_trigger_
        array_obj_ref_486_active_x_x2118_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_active_ 
          signal array_obj_ref_486_active_x_x2118_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_486_active_x_x2118_predecessors(0) <= array_obj_ref_486_trigger_x_x2117_symbol;
          array_obj_ref_486_active_x_x2118_predecessors(1) <= array_obj_ref_486_root_address_calculated_2120_symbol;
          array_obj_ref_486_active_x_x2118_join: join -- 
            port map( -- 
              preds => array_obj_ref_486_active_x_x2118_predecessors,
              symbol_out => array_obj_ref_486_active_x_x2118_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_active_
        array_obj_ref_486_base_address_calculated_2119_symbol <= assign_stmt_482_completed_x_x2085_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_address_calculated
        array_obj_ref_486_root_address_calculated_2120_symbol <= array_obj_ref_486_base_plus_offset_2128_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_root_address_calculated
        array_obj_ref_486_base_address_resized_2121_symbol <= array_obj_ref_486_base_addr_resize_2122_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_address_resized
        array_obj_ref_486_base_addr_resize_2122: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize 
          signal array_obj_ref_486_base_addr_resize_2122_start: Boolean;
          signal Xentry_2123_symbol: Boolean;
          signal Xexit_2124_symbol: Boolean;
          signal base_resize_req_2125_symbol : Boolean;
          signal base_resize_ack_2126_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_486_base_addr_resize_2122_start <= array_obj_ref_486_base_address_calculated_2119_symbol; -- control passed to block
          Xentry_2123_symbol  <= array_obj_ref_486_base_addr_resize_2122_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/$entry
          base_resize_req_2125_symbol <= Xentry_2123_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/base_resize_req
          array_obj_ref_486_base_resize_req_0 <= base_resize_req_2125_symbol; -- link to DP
          base_resize_ack_2126_symbol <= array_obj_ref_486_base_resize_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/base_resize_ack
          Xexit_2124_symbol <= base_resize_ack_2126_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize/$exit
          array_obj_ref_486_base_addr_resize_2122_symbol <= Xexit_2124_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_addr_resize
        array_obj_ref_486_base_plus_offset_trigger_2127_symbol <= array_obj_ref_486_base_address_resized_2121_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset_trigger
        array_obj_ref_486_base_plus_offset_2128: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset 
          signal array_obj_ref_486_base_plus_offset_2128_start: Boolean;
          signal Xentry_2129_symbol: Boolean;
          signal Xexit_2130_symbol: Boolean;
          signal plus_base_rr_2131_symbol : Boolean;
          signal plus_base_ra_2132_symbol : Boolean;
          signal plus_base_cr_2133_symbol : Boolean;
          signal plus_base_ca_2134_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_486_base_plus_offset_2128_start <= array_obj_ref_486_base_plus_offset_trigger_2127_symbol; -- control passed to block
          Xentry_2129_symbol  <= array_obj_ref_486_base_plus_offset_2128_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/$entry
          plus_base_rr_2131_symbol <= Xentry_2129_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_rr
          array_obj_ref_486_root_address_inst_req_0 <= plus_base_rr_2131_symbol; -- link to DP
          plus_base_ra_2132_symbol <= array_obj_ref_486_root_address_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_ra
          plus_base_cr_2133_symbol <= plus_base_ra_2132_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_cr
          array_obj_ref_486_root_address_inst_req_1 <= plus_base_cr_2133_symbol; -- link to DP
          plus_base_ca_2134_symbol <= array_obj_ref_486_root_address_inst_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/plus_base_ca
          Xexit_2130_symbol <= plus_base_ca_2134_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset/$exit
          array_obj_ref_486_base_plus_offset_2128_symbol <= Xexit_2130_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_base_plus_offset
        array_obj_ref_486_complete_2135: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete 
          signal array_obj_ref_486_complete_2135_start: Boolean;
          signal Xentry_2136_symbol: Boolean;
          signal Xexit_2137_symbol: Boolean;
          signal final_reg_req_2138_symbol : Boolean;
          signal final_reg_ack_2139_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_486_complete_2135_start <= array_obj_ref_486_active_x_x2118_symbol; -- control passed to block
          Xentry_2136_symbol  <= array_obj_ref_486_complete_2135_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/$entry
          final_reg_req_2138_symbol <= Xentry_2136_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/final_reg_req
          array_obj_ref_486_final_reg_req_0 <= final_reg_req_2138_symbol; -- link to DP
          final_reg_ack_2139_symbol <= array_obj_ref_486_final_reg_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/final_reg_ack
          Xexit_2137_symbol <= final_reg_ack_2139_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete/$exit
          array_obj_ref_486_complete_2135_symbol <= Xexit_2137_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/array_obj_ref_486_complete
        assign_stmt_491_active_x_x2140_symbol <= simple_obj_ref_490_complete_2142_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_491_active_
        assign_stmt_491_completed_x_x2141_symbol <= ptr_deref_489_complete_2178_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_491_completed_
        simple_obj_ref_490_complete_2142_symbol <= assign_stmt_478_completed_x_x2054_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_490_complete
        ptr_deref_489_trigger_x_x2143_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_trigger_ 
          signal ptr_deref_489_trigger_x_x2143_predecessors: BooleanArray(2 downto 0);
          -- 
        begin -- 
          ptr_deref_489_trigger_x_x2143_predecessors(0) <= ptr_deref_489_word_address_calculated_2148_symbol;
          ptr_deref_489_trigger_x_x2143_predecessors(1) <= ptr_deref_489_base_address_calculated_2145_symbol;
          ptr_deref_489_trigger_x_x2143_predecessors(2) <= assign_stmt_491_active_x_x2140_symbol;
          ptr_deref_489_trigger_x_x2143_join: join -- 
            port map( -- 
              preds => ptr_deref_489_trigger_x_x2143_predecessors,
              symbol_out => ptr_deref_489_trigger_x_x2143_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_trigger_
        ptr_deref_489_active_x_x2144_symbol <= ptr_deref_489_request_2165_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_active_
        ptr_deref_489_base_address_calculated_2145_symbol <= simple_obj_ref_488_complete_2146_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_address_calculated
        simple_obj_ref_488_complete_2146_symbol <= assign_stmt_487_completed_x_x2116_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_488_complete
        ptr_deref_489_root_address_calculated_2147_symbol <= ptr_deref_489_base_plus_offset_2155_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_root_address_calculated
        ptr_deref_489_word_address_calculated_2148_symbol <= ptr_deref_489_word_addrgen_2160_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_address_calculated
        ptr_deref_489_base_address_resized_2149_symbol <= ptr_deref_489_base_addr_resize_2150_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_address_resized
        ptr_deref_489_base_addr_resize_2150: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize 
          signal ptr_deref_489_base_addr_resize_2150_start: Boolean;
          signal Xentry_2151_symbol: Boolean;
          signal Xexit_2152_symbol: Boolean;
          signal base_resize_req_2153_symbol : Boolean;
          signal base_resize_ack_2154_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_base_addr_resize_2150_start <= ptr_deref_489_base_address_calculated_2145_symbol; -- control passed to block
          Xentry_2151_symbol  <= ptr_deref_489_base_addr_resize_2150_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/$entry
          base_resize_req_2153_symbol <= Xentry_2151_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/base_resize_req
          ptr_deref_489_base_resize_req_0 <= base_resize_req_2153_symbol; -- link to DP
          base_resize_ack_2154_symbol <= ptr_deref_489_base_resize_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/base_resize_ack
          Xexit_2152_symbol <= base_resize_ack_2154_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize/$exit
          ptr_deref_489_base_addr_resize_2150_symbol <= Xexit_2152_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_addr_resize
        ptr_deref_489_base_plus_offset_2155: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset 
          signal ptr_deref_489_base_plus_offset_2155_start: Boolean;
          signal Xentry_2156_symbol: Boolean;
          signal Xexit_2157_symbol: Boolean;
          signal sum_rename_req_2158_symbol : Boolean;
          signal sum_rename_ack_2159_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_base_plus_offset_2155_start <= ptr_deref_489_base_address_resized_2149_symbol; -- control passed to block
          Xentry_2156_symbol  <= ptr_deref_489_base_plus_offset_2155_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/$entry
          sum_rename_req_2158_symbol <= Xentry_2156_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/sum_rename_req
          ptr_deref_489_root_address_inst_req_0 <= sum_rename_req_2158_symbol; -- link to DP
          sum_rename_ack_2159_symbol <= ptr_deref_489_root_address_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/sum_rename_ack
          Xexit_2157_symbol <= sum_rename_ack_2159_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset/$exit
          ptr_deref_489_base_plus_offset_2155_symbol <= Xexit_2157_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_base_plus_offset
        ptr_deref_489_word_addrgen_2160: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen 
          signal ptr_deref_489_word_addrgen_2160_start: Boolean;
          signal Xentry_2161_symbol: Boolean;
          signal Xexit_2162_symbol: Boolean;
          signal root_rename_req_2163_symbol : Boolean;
          signal root_rename_ack_2164_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_word_addrgen_2160_start <= ptr_deref_489_root_address_calculated_2147_symbol; -- control passed to block
          Xentry_2161_symbol  <= ptr_deref_489_word_addrgen_2160_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/$entry
          root_rename_req_2163_symbol <= Xentry_2161_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/root_rename_req
          ptr_deref_489_addr_0_req_0 <= root_rename_req_2163_symbol; -- link to DP
          root_rename_ack_2164_symbol <= ptr_deref_489_addr_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/root_rename_ack
          Xexit_2162_symbol <= root_rename_ack_2164_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen/$exit
          ptr_deref_489_word_addrgen_2160_symbol <= Xexit_2162_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_word_addrgen
        ptr_deref_489_request_2165: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request 
          signal ptr_deref_489_request_2165_start: Boolean;
          signal Xentry_2166_symbol: Boolean;
          signal Xexit_2167_symbol: Boolean;
          signal split_req_2168_symbol : Boolean;
          signal split_ack_2169_symbol : Boolean;
          signal word_access_2170_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_request_2165_start <= ptr_deref_489_trigger_x_x2143_symbol; -- control passed to block
          Xentry_2166_symbol  <= ptr_deref_489_request_2165_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/$entry
          split_req_2168_symbol <= Xentry_2166_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/split_req
          ptr_deref_489_gather_scatter_req_0 <= split_req_2168_symbol; -- link to DP
          split_ack_2169_symbol <= ptr_deref_489_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/split_ack
          word_access_2170: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access 
            signal word_access_2170_start: Boolean;
            signal Xentry_2171_symbol: Boolean;
            signal Xexit_2172_symbol: Boolean;
            signal word_access_0_2173_symbol : Boolean;
            -- 
          begin -- 
            word_access_2170_start <= split_ack_2169_symbol; -- control passed to block
            Xentry_2171_symbol  <= word_access_2170_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/$entry
            word_access_0_2173: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0 
              signal word_access_0_2173_start: Boolean;
              signal Xentry_2174_symbol: Boolean;
              signal Xexit_2175_symbol: Boolean;
              signal rr_2176_symbol : Boolean;
              signal ra_2177_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2173_start <= Xentry_2171_symbol; -- control passed to block
              Xentry_2174_symbol  <= word_access_0_2173_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/$entry
              rr_2176_symbol <= Xentry_2174_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/rr
              ptr_deref_489_store_0_req_0 <= rr_2176_symbol; -- link to DP
              ra_2177_symbol <= ptr_deref_489_store_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/ra
              Xexit_2175_symbol <= ra_2177_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0/$exit
              word_access_0_2173_symbol <= Xexit_2175_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/word_access_0
            Xexit_2172_symbol <= word_access_0_2173_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access/$exit
            word_access_2170_symbol <= Xexit_2172_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/word_access
          Xexit_2167_symbol <= word_access_2170_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request/$exit
          ptr_deref_489_request_2165_symbol <= Xexit_2167_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_request
        ptr_deref_489_complete_2178: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete 
          signal ptr_deref_489_complete_2178_start: Boolean;
          signal Xentry_2179_symbol: Boolean;
          signal Xexit_2180_symbol: Boolean;
          signal word_access_2181_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_489_complete_2178_start <= ptr_deref_489_active_x_x2144_symbol; -- control passed to block
          Xentry_2179_symbol  <= ptr_deref_489_complete_2178_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/$entry
          word_access_2181: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access 
            signal word_access_2181_start: Boolean;
            signal Xentry_2182_symbol: Boolean;
            signal Xexit_2183_symbol: Boolean;
            signal word_access_0_2184_symbol : Boolean;
            -- 
          begin -- 
            word_access_2181_start <= Xentry_2179_symbol; -- control passed to block
            Xentry_2182_symbol  <= word_access_2181_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/$entry
            word_access_0_2184: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0 
              signal word_access_0_2184_start: Boolean;
              signal Xentry_2185_symbol: Boolean;
              signal Xexit_2186_symbol: Boolean;
              signal cr_2187_symbol : Boolean;
              signal ca_2188_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2184_start <= Xentry_2182_symbol; -- control passed to block
              Xentry_2185_symbol  <= word_access_0_2184_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/$entry
              cr_2187_symbol <= Xentry_2185_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/cr
              ptr_deref_489_store_0_req_1 <= cr_2187_symbol; -- link to DP
              ca_2188_symbol <= ptr_deref_489_store_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/ca
              Xexit_2186_symbol <= ca_2188_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0/$exit
              word_access_0_2184_symbol <= Xexit_2186_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/word_access_0
            Xexit_2183_symbol <= word_access_0_2184_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access/$exit
            word_access_2181_symbol <= Xexit_2183_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/word_access
          Xexit_2180_symbol <= word_access_2181_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete/$exit
          ptr_deref_489_complete_2178_symbol <= Xexit_2180_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_489_complete
        assign_stmt_495_active_x_x2189_symbol <= ptr_deref_494_complete_2207_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_495_active_
        assign_stmt_495_completed_x_x2190_symbol <= assign_stmt_495_active_x_x2189_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_495_completed_
        ptr_deref_494_trigger_x_x2191_symbol <= ptr_deref_494_word_address_calculated_2195_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_trigger_
        ptr_deref_494_active_x_x2192_symbol <= ptr_deref_494_request_2196_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_active_
        ptr_deref_494_base_address_calculated_2193_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_base_address_calculated
        ptr_deref_494_root_address_calculated_2194_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_root_address_calculated
        ptr_deref_494_word_address_calculated_2195_symbol <= ptr_deref_494_root_address_calculated_2194_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_word_address_calculated
        ptr_deref_494_request_2196: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request 
          signal ptr_deref_494_request_2196_start: Boolean;
          signal Xentry_2197_symbol: Boolean;
          signal Xexit_2198_symbol: Boolean;
          signal word_access_2199_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_494_request_2196_start <= ptr_deref_494_trigger_x_x2191_symbol; -- control passed to block
          Xentry_2197_symbol  <= ptr_deref_494_request_2196_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/$entry
          word_access_2199: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access 
            signal word_access_2199_start: Boolean;
            signal Xentry_2200_symbol: Boolean;
            signal Xexit_2201_symbol: Boolean;
            signal word_access_0_2202_symbol : Boolean;
            -- 
          begin -- 
            word_access_2199_start <= Xentry_2197_symbol; -- control passed to block
            Xentry_2200_symbol  <= word_access_2199_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/$entry
            word_access_0_2202: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0 
              signal word_access_0_2202_start: Boolean;
              signal Xentry_2203_symbol: Boolean;
              signal Xexit_2204_symbol: Boolean;
              signal rr_2205_symbol : Boolean;
              signal ra_2206_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2202_start <= Xentry_2200_symbol; -- control passed to block
              Xentry_2203_symbol  <= word_access_0_2202_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/$entry
              rr_2205_symbol <= Xentry_2203_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/rr
              ptr_deref_494_load_0_req_0 <= rr_2205_symbol; -- link to DP
              ra_2206_symbol <= ptr_deref_494_load_0_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/ra
              Xexit_2204_symbol <= ra_2206_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0/$exit
              word_access_0_2202_symbol <= Xexit_2204_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/word_access_0
            Xexit_2201_symbol <= word_access_0_2202_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access/$exit
            word_access_2199_symbol <= Xexit_2201_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/word_access
          Xexit_2198_symbol <= word_access_2199_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request/$exit
          ptr_deref_494_request_2196_symbol <= Xexit_2198_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_request
        ptr_deref_494_complete_2207: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete 
          signal ptr_deref_494_complete_2207_start: Boolean;
          signal Xentry_2208_symbol: Boolean;
          signal Xexit_2209_symbol: Boolean;
          signal word_access_2210_symbol : Boolean;
          signal merge_req_2218_symbol : Boolean;
          signal merge_ack_2219_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_494_complete_2207_start <= ptr_deref_494_active_x_x2192_symbol; -- control passed to block
          Xentry_2208_symbol  <= ptr_deref_494_complete_2207_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/$entry
          word_access_2210: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access 
            signal word_access_2210_start: Boolean;
            signal Xentry_2211_symbol: Boolean;
            signal Xexit_2212_symbol: Boolean;
            signal word_access_0_2213_symbol : Boolean;
            -- 
          begin -- 
            word_access_2210_start <= Xentry_2208_symbol; -- control passed to block
            Xentry_2211_symbol  <= word_access_2210_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/$entry
            word_access_0_2213: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0 
              signal word_access_0_2213_start: Boolean;
              signal Xentry_2214_symbol: Boolean;
              signal Xexit_2215_symbol: Boolean;
              signal cr_2216_symbol : Boolean;
              signal ca_2217_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2213_start <= Xentry_2211_symbol; -- control passed to block
              Xentry_2214_symbol  <= word_access_0_2213_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/$entry
              cr_2216_symbol <= Xentry_2214_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/cr
              ptr_deref_494_load_0_req_1 <= cr_2216_symbol; -- link to DP
              ca_2217_symbol <= ptr_deref_494_load_0_ack_1; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/ca
              Xexit_2215_symbol <= ca_2217_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0/$exit
              word_access_0_2213_symbol <= Xexit_2215_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/word_access_0
            Xexit_2212_symbol <= word_access_0_2213_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access/$exit
            word_access_2210_symbol <= Xexit_2212_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/word_access
          merge_req_2218_symbol <= word_access_2210_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/merge_req
          ptr_deref_494_gather_scatter_req_0 <= merge_req_2218_symbol; -- link to DP
          merge_ack_2219_symbol <= ptr_deref_494_gather_scatter_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/merge_ack
          Xexit_2209_symbol <= merge_ack_2219_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete/$exit
          ptr_deref_494_complete_2207_symbol <= Xexit_2209_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/ptr_deref_494_complete
        assign_stmt_499_active_x_x2220_symbol <= type_cast_498_complete_2225_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_499_active_
        assign_stmt_499_completed_x_x2221_symbol <= assign_stmt_499_active_x_x2220_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/assign_stmt_499_completed_
        type_cast_498_active_x_x2222_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_active_ 
          signal type_cast_498_active_x_x2222_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_498_active_x_x2222_predecessors(0) <= type_cast_498_trigger_x_x2223_symbol;
          type_cast_498_active_x_x2222_predecessors(1) <= simple_obj_ref_497_complete_2224_symbol;
          type_cast_498_active_x_x2222_join: join -- 
            port map( -- 
              preds => type_cast_498_active_x_x2222_predecessors,
              symbol_out => type_cast_498_active_x_x2222_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_active_
        type_cast_498_trigger_x_x2223_symbol <= Xentry_2019_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_trigger_
        simple_obj_ref_497_complete_2224_symbol <= assign_stmt_495_completed_x_x2190_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/simple_obj_ref_497_complete
        type_cast_498_complete_2225: Block -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete 
          signal type_cast_498_complete_2225_start: Boolean;
          signal Xentry_2226_symbol: Boolean;
          signal Xexit_2227_symbol: Boolean;
          signal req_2228_symbol : Boolean;
          signal ack_2229_symbol : Boolean;
          -- 
        begin -- 
          type_cast_498_complete_2225_start <= type_cast_498_active_x_x2222_symbol; -- control passed to block
          Xentry_2226_symbol  <= type_cast_498_complete_2225_start; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/$entry
          req_2228_symbol <= Xentry_2226_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/req
          type_cast_498_inst_req_0 <= req_2228_symbol; -- link to DP
          ack_2229_symbol <= type_cast_498_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/ack
          Xexit_2227_symbol <= ack_2229_symbol; -- transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete/$exit
          type_cast_498_complete_2225_symbol <= Xexit_2227_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/type_cast_498_complete
        Xexit_2020_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/$exit 
          signal Xexit_2020_predecessors: BooleanArray(6 downto 0);
          -- 
        begin -- 
          Xexit_2020_predecessors(0) <= assign_stmt_474_completed_x_x2022_symbol;
          Xexit_2020_predecessors(1) <= ptr_deref_472_base_address_calculated_2026_symbol;
          Xexit_2020_predecessors(2) <= ptr_deref_477_base_address_calculated_2057_symbol;
          Xexit_2020_predecessors(3) <= ptr_deref_481_base_address_calculated_2088_symbol;
          Xexit_2020_predecessors(4) <= assign_stmt_491_completed_x_x2141_symbol;
          Xexit_2020_predecessors(5) <= ptr_deref_494_base_address_calculated_2193_symbol;
          Xexit_2020_predecessors(6) <= assign_stmt_499_completed_x_x2221_symbol;
          Xexit_2020_join: join -- 
            port map( -- 
              preds => Xexit_2020_predecessors,
              symbol_out => Xexit_2020_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504/$exit
        assign_stmt_474_to_assign_stmt_504_2018_symbol <= Xexit_2020_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_474_to_assign_stmt_504
      assign_stmt_508_2230: Block -- branch_block_stmt_405/assign_stmt_508 
        signal assign_stmt_508_2230_start: Boolean;
        signal Xentry_2231_symbol: Boolean;
        signal Xexit_2232_symbol: Boolean;
        signal assign_stmt_508_active_x_x2233_symbol : Boolean;
        signal assign_stmt_508_completed_x_x2234_symbol : Boolean;
        signal type_cast_507_active_x_x2235_symbol : Boolean;
        signal type_cast_507_trigger_x_x2236_symbol : Boolean;
        signal simple_obj_ref_506_complete_2237_symbol : Boolean;
        signal type_cast_507_complete_2238_symbol : Boolean;
        signal simple_obj_ref_505_trigger_x_x2243_symbol : Boolean;
        signal simple_obj_ref_505_complete_2244_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_508_2230_start <= assign_stmt_508_x_xentry_x_xx_x1842_symbol; -- control passed to block
        Xentry_2231_symbol  <= assign_stmt_508_2230_start; -- transition branch_block_stmt_405/assign_stmt_508/$entry
        assign_stmt_508_active_x_x2233_symbol <= type_cast_507_complete_2238_symbol; -- transition branch_block_stmt_405/assign_stmt_508/assign_stmt_508_active_
        assign_stmt_508_completed_x_x2234_symbol <= simple_obj_ref_505_complete_2244_symbol; -- transition branch_block_stmt_405/assign_stmt_508/assign_stmt_508_completed_
        type_cast_507_active_x_x2235_block : Block -- non-trivial join transition branch_block_stmt_405/assign_stmt_508/type_cast_507_active_ 
          signal type_cast_507_active_x_x2235_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_507_active_x_x2235_predecessors(0) <= type_cast_507_trigger_x_x2236_symbol;
          type_cast_507_active_x_x2235_predecessors(1) <= simple_obj_ref_506_complete_2237_symbol;
          type_cast_507_active_x_x2235_join: join -- 
            port map( -- 
              preds => type_cast_507_active_x_x2235_predecessors,
              symbol_out => type_cast_507_active_x_x2235_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_405/assign_stmt_508/type_cast_507_active_
        type_cast_507_trigger_x_x2236_symbol <= Xentry_2231_symbol; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_trigger_
        simple_obj_ref_506_complete_2237_symbol <= Xentry_2231_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_506_complete
        type_cast_507_complete_2238: Block -- branch_block_stmt_405/assign_stmt_508/type_cast_507_complete 
          signal type_cast_507_complete_2238_start: Boolean;
          signal Xentry_2239_symbol: Boolean;
          signal Xexit_2240_symbol: Boolean;
          signal req_2241_symbol : Boolean;
          signal ack_2242_symbol : Boolean;
          -- 
        begin -- 
          type_cast_507_complete_2238_start <= type_cast_507_active_x_x2235_symbol; -- control passed to block
          Xentry_2239_symbol  <= type_cast_507_complete_2238_start; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/$entry
          req_2241_symbol <= Xentry_2239_symbol; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/req
          type_cast_507_inst_req_0 <= req_2241_symbol; -- link to DP
          ack_2242_symbol <= type_cast_507_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/ack
          Xexit_2240_symbol <= ack_2242_symbol; -- transition branch_block_stmt_405/assign_stmt_508/type_cast_507_complete/$exit
          type_cast_507_complete_2238_symbol <= Xexit_2240_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_508/type_cast_507_complete
        simple_obj_ref_505_trigger_x_x2243_symbol <= assign_stmt_508_active_x_x2233_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_trigger_
        simple_obj_ref_505_complete_2244: Block -- branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete 
          signal simple_obj_ref_505_complete_2244_start: Boolean;
          signal Xentry_2245_symbol: Boolean;
          signal Xexit_2246_symbol: Boolean;
          signal pipe_wreq_2247_symbol : Boolean;
          signal pipe_wack_2248_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_505_complete_2244_start <= simple_obj_ref_505_trigger_x_x2243_symbol; -- control passed to block
          Xentry_2245_symbol  <= simple_obj_ref_505_complete_2244_start; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/$entry
          pipe_wreq_2247_symbol <= Xentry_2245_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/pipe_wreq
          simple_obj_ref_505_inst_req_0 <= pipe_wreq_2247_symbol; -- link to DP
          pipe_wack_2248_symbol <= simple_obj_ref_505_inst_ack_0; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/pipe_wack
          Xexit_2246_symbol <= pipe_wack_2248_symbol; -- transition branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete/$exit
          simple_obj_ref_505_complete_2244_symbol <= Xexit_2246_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_405/assign_stmt_508/simple_obj_ref_505_complete
        Xexit_2232_symbol <= assign_stmt_508_completed_x_x2234_symbol; -- transition branch_block_stmt_405/assign_stmt_508/$exit
        assign_stmt_508_2230_symbol <= Xexit_2232_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/assign_stmt_508
      bb_0_bb_1_PhiReq_2249: Block -- branch_block_stmt_405/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_2249_start: Boolean;
        signal Xentry_2250_symbol: Boolean;
        signal Xexit_2251_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_2249_start <= bb_0_bb_1_1820_symbol; -- control passed to block
        Xentry_2250_symbol  <= bb_0_bb_1_PhiReq_2249_start; -- transition branch_block_stmt_405/bb_0_bb_1_PhiReq/$entry
        Xexit_2251_symbol <= Xentry_2250_symbol; -- transition branch_block_stmt_405/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_2249_symbol <= Xexit_2251_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_0_bb_1_PhiReq
      bb_1_bb_1_PhiReq_2252: Block -- branch_block_stmt_405/bb_1_bb_1_PhiReq 
        signal bb_1_bb_1_PhiReq_2252_start: Boolean;
        signal Xentry_2253_symbol: Boolean;
        signal Xexit_2254_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_1_PhiReq_2252_start <= bb_1_bb_1_1996_symbol; -- control passed to block
        Xentry_2253_symbol  <= bb_1_bb_1_PhiReq_2252_start; -- transition branch_block_stmt_405/bb_1_bb_1_PhiReq/$entry
        Xexit_2254_symbol <= Xentry_2253_symbol; -- transition branch_block_stmt_405/bb_1_bb_1_PhiReq/$exit
        bb_1_bb_1_PhiReq_2252_symbol <= Xexit_2254_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_1_bb_1_PhiReq
      bb_2_bb_1_PhiReq_2255: Block -- branch_block_stmt_405/bb_2_bb_1_PhiReq 
        signal bb_2_bb_1_PhiReq_2255_start: Boolean;
        signal Xentry_2256_symbol: Boolean;
        signal Xexit_2257_symbol: Boolean;
        -- 
      begin -- 
        bb_2_bb_1_PhiReq_2255_start <= bb_2_bb_1_1844_symbol; -- control passed to block
        Xentry_2256_symbol  <= bb_2_bb_1_PhiReq_2255_start; -- transition branch_block_stmt_405/bb_2_bb_1_PhiReq/$entry
        Xexit_2257_symbol <= Xentry_2256_symbol; -- transition branch_block_stmt_405/bb_2_bb_1_PhiReq/$exit
        bb_2_bb_1_PhiReq_2255_symbol <= Xexit_2257_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_2_bb_1_PhiReq
      merge_stmt_417_PhiReqMerge_2258_symbol  <=  bb_0_bb_1_PhiReq_2249_symbol or bb_1_bb_1_PhiReq_2252_symbol or bb_2_bb_1_PhiReq_2255_symbol; -- place branch_block_stmt_405/merge_stmt_417_PhiReqMerge (optimized away) 
      merge_stmt_417_PhiAck_2259: Block -- branch_block_stmt_405/merge_stmt_417_PhiAck 
        signal merge_stmt_417_PhiAck_2259_start: Boolean;
        signal Xentry_2260_symbol: Boolean;
        signal Xexit_2261_symbol: Boolean;
        signal dummy_2262_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_417_PhiAck_2259_start <= merge_stmt_417_PhiReqMerge_2258_symbol; -- control passed to block
        Xentry_2260_symbol  <= merge_stmt_417_PhiAck_2259_start; -- transition branch_block_stmt_405/merge_stmt_417_PhiAck/$entry
        dummy_2262_symbol <= Xentry_2260_symbol; -- transition branch_block_stmt_405/merge_stmt_417_PhiAck/dummy
        Xexit_2261_symbol <= dummy_2262_symbol; -- transition branch_block_stmt_405/merge_stmt_417_PhiAck/$exit
        merge_stmt_417_PhiAck_2259_symbol <= Xexit_2261_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/merge_stmt_417_PhiAck
      merge_stmt_461_dead_link_2263: Block -- branch_block_stmt_405/merge_stmt_461_dead_link 
        signal merge_stmt_461_dead_link_2263_start: Boolean;
        signal Xentry_2264_symbol: Boolean;
        signal Xexit_2265_symbol: Boolean;
        signal dead_transition_2266_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_461_dead_link_2263_start <= merge_stmt_461_x_xentry_x_xx_x1834_symbol; -- control passed to block
        Xentry_2264_symbol  <= merge_stmt_461_dead_link_2263_start; -- transition branch_block_stmt_405/merge_stmt_461_dead_link/$entry
        dead_transition_2266_symbol <= false;
        Xexit_2265_symbol <= dead_transition_2266_symbol; -- transition branch_block_stmt_405/merge_stmt_461_dead_link/$exit
        merge_stmt_461_dead_link_2263_symbol <= Xexit_2265_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/merge_stmt_461_dead_link
      bb_1_bb_2_PhiReq_2267: Block -- branch_block_stmt_405/bb_1_bb_2_PhiReq 
        signal bb_1_bb_2_PhiReq_2267_start: Boolean;
        signal Xentry_2268_symbol: Boolean;
        signal Xexit_2269_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_2_PhiReq_2267_start <= bb_1_bb_2_1995_symbol; -- control passed to block
        Xentry_2268_symbol  <= bb_1_bb_2_PhiReq_2267_start; -- transition branch_block_stmt_405/bb_1_bb_2_PhiReq/$entry
        Xexit_2269_symbol <= Xentry_2268_symbol; -- transition branch_block_stmt_405/bb_1_bb_2_PhiReq/$exit
        bb_1_bb_2_PhiReq_2267_symbol <= Xexit_2269_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/bb_1_bb_2_PhiReq
      merge_stmt_461_PhiReqMerge_2270_symbol  <=  bb_1_bb_2_PhiReq_2267_symbol; -- place branch_block_stmt_405/merge_stmt_461_PhiReqMerge (optimized away) 
      merge_stmt_461_PhiAck_2271: Block -- branch_block_stmt_405/merge_stmt_461_PhiAck 
        signal merge_stmt_461_PhiAck_2271_start: Boolean;
        signal Xentry_2272_symbol: Boolean;
        signal Xexit_2273_symbol: Boolean;
        signal dummy_2274_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_461_PhiAck_2271_start <= merge_stmt_461_PhiReqMerge_2270_symbol; -- control passed to block
        Xentry_2272_symbol  <= merge_stmt_461_PhiAck_2271_start; -- transition branch_block_stmt_405/merge_stmt_461_PhiAck/$entry
        dummy_2274_symbol <= Xentry_2272_symbol; -- transition branch_block_stmt_405/merge_stmt_461_PhiAck/dummy
        Xexit_2273_symbol <= dummy_2274_symbol; -- transition branch_block_stmt_405/merge_stmt_461_PhiAck/$exit
        merge_stmt_461_PhiAck_2271_symbol <= Xexit_2273_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_405/merge_stmt_461_PhiAck
      Xexit_1815_symbol <= branch_block_stmt_405_x_xexit_x_xx_x1817_symbol; -- transition branch_block_stmt_405/$exit
      branch_block_stmt_405_1813_symbol <= Xexit_1815_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_405
    Xexit_1812_symbol <= branch_block_stmt_405_1813_symbol; -- transition $exit
    fin  <=  '1' when Xexit_1812_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_486_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_486_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_486_root_address : std_logic_vector(2 downto 0);
    signal iNsTr_10_466 : std_logic_vector(31 downto 0);
    signal iNsTr_11_470 : std_logic_vector(31 downto 0);
    signal iNsTr_13_478 : std_logic_vector(31 downto 0);
    signal iNsTr_14_482 : std_logic_vector(31 downto 0);
    signal iNsTr_15_487 : std_logic_vector(31 downto 0);
    signal iNsTr_17_495 : std_logic_vector(31 downto 0);
    signal iNsTr_18_499 : std_logic_vector(31 downto 0);
    signal iNsTr_19_504 : std_logic_vector(31 downto 0);
    signal iNsTr_1_422 : std_logic_vector(31 downto 0);
    signal iNsTr_3_431 : std_logic_vector(31 downto 0);
    signal iNsTr_4_435 : std_logic_vector(31 downto 0);
    signal iNsTr_5_439 : std_logic_vector(31 downto 0);
    signal iNsTr_7_447 : std_logic_vector(31 downto 0);
    signal iNsTr_8_454 : std_logic_vector(0 downto 0);
    signal lptr_411 : std_logic_vector(31 downto 0);
    signal nval_415 : std_logic_vector(31 downto 0);
    signal ptr_deref_441_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_441_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_441_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_446_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_446_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_472_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_472_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_472_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_477_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_477_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_481_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_481_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_489_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_489_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_489_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_489_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_489_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_489_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_494_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_494_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_433_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_468_wire : std_logic_vector(31 downto 0);
    signal type_cast_425_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_450_wire : std_logic_vector(31 downto 0);
    signal type_cast_452_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_507_wire : std_logic_vector(31 downto 0);
    signal xxinput_modulexxbodyxxlptr_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxinput_modulexxbodyxxnval_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_486_final_offset <= "001";
    iNsTr_10_466 <= "00000000000000000000000000000000";
    iNsTr_19_504 <= "00000000000000000000000000000000";
    iNsTr_1_422 <= "00000000000000000000000000000000";
    iNsTr_3_431 <= "00000000000000000000000000000000";
    lptr_411 <= "00000000000000000000000000000000";
    nval_415 <= "00000000000000000000000000000000";
    ptr_deref_441_word_address_0 <= "0";
    ptr_deref_446_word_address_0 <= "0";
    ptr_deref_472_word_address_0 <= "0";
    ptr_deref_477_word_address_0 <= "0";
    ptr_deref_481_word_address_0 <= "0";
    ptr_deref_489_word_offset_0 <= "000";
    ptr_deref_494_word_address_0 <= "0";
    type_cast_425_wire_constant <= "00000010";
    type_cast_452_wire_constant <= "11111111111111111111111111111111";
    xxinput_modulexxbodyxxlptr_alloc_base_address <= "0";
    xxinput_modulexxbodyxxnval_alloc_base_address <= "0";
    array_obj_ref_486_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_14_482, dout => array_obj_ref_486_resized_base_address, req => array_obj_ref_486_base_resize_req_0, ack => array_obj_ref_486_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_486_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_486_root_address, dout => iNsTr_15_487, req => array_obj_ref_486_final_reg_req_0, ack => array_obj_ref_486_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_489_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_15_487, dout => ptr_deref_489_resized_base_address, req => ptr_deref_489_base_resize_req_0, ack => ptr_deref_489_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_434_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_433_wire, dout => iNsTr_4_435, req => type_cast_434_inst_req_0, ack => type_cast_434_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_438_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_4_435, dout => iNsTr_5_439, req => type_cast_438_inst_req_0, ack => type_cast_438_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_450_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_7_447, dout => type_cast_450_wire, req => type_cast_450_inst_req_0, ack => type_cast_450_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_469_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_468_wire, dout => iNsTr_11_470, req => type_cast_469_inst_req_0, ack => type_cast_469_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_498_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_17_495, dout => iNsTr_18_499, req => type_cast_498_inst_req_0, ack => type_cast_498_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_507_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_18_499, dout => type_cast_507_wire, req => type_cast_507_inst_req_0, ack => type_cast_507_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_441_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_441_gather_scatter_ack_0 <= ptr_deref_441_gather_scatter_req_0;
      aggregated_sig <= iNsTr_5_439;
      ptr_deref_441_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_446_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_446_gather_scatter_ack_0 <= ptr_deref_446_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_446_data_0;
      iNsTr_7_447 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_472_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_472_gather_scatter_ack_0 <= ptr_deref_472_gather_scatter_req_0;
      aggregated_sig <= iNsTr_11_470;
      ptr_deref_472_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_477_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_477_gather_scatter_ack_0 <= ptr_deref_477_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_477_data_0;
      iNsTr_13_478 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_481_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_481_gather_scatter_ack_0 <= ptr_deref_481_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_481_data_0;
      iNsTr_14_482 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_489_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_489_addr_0_ack_0 <= ptr_deref_489_addr_0_req_0;
      aggregated_sig <= ptr_deref_489_root_address;
      ptr_deref_489_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_489_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_489_gather_scatter_ack_0 <= ptr_deref_489_gather_scatter_req_0;
      aggregated_sig <= iNsTr_13_478;
      ptr_deref_489_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_489_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_489_root_address_inst_ack_0 <= ptr_deref_489_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_489_resized_base_address;
      ptr_deref_489_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_494_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_494_gather_scatter_ack_0 <= ptr_deref_494_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_494_data_0;
      iNsTr_17_495 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_455_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_8_454;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_455_branch_req_0,
          ack0 => if_stmt_455_branch_ack_0,
          ack1 => if_stmt_455_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_486_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_486_resized_base_address;
      array_obj_ref_486_root_address <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_486_root_address_inst_req_0,
          ackL => array_obj_ref_486_root_address_inst_ack_0,
          reqR => array_obj_ref_486_root_address_inst_req_1,
          ackR => array_obj_ref_486_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_453_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_450_wire;
      iNsTr_8_454 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_453_inst_req_0,
          ackL => binary_453_inst_ack_0,
          reqR => binary_453_inst_req_1,
          ackR => binary_453_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared load operator group (0) : ptr_deref_446_load_0 ptr_deref_481_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_446_load_0_req_0;
      reqL(0) <= ptr_deref_481_load_0_req_0;
      ptr_deref_446_load_0_ack_0 <= ackL(1);
      ptr_deref_481_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_446_load_0_req_1;
      reqR(0) <= ptr_deref_481_load_0_req_1;
      ptr_deref_446_load_0_ack_1 <= ackR(1);
      ptr_deref_481_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_446_word_address_0 & ptr_deref_481_word_address_0;
      ptr_deref_446_data_0 <= data_out(63 downto 32);
      ptr_deref_481_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_15_lr_req(1),
          mack => memory_space_15_lr_ack(1),
          maddr => memory_space_15_lr_addr(1 downto 1),
          mtag => memory_space_15_lr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_15_lc_req(1),
          mack => memory_space_15_lc_ack(1),
          mdata => memory_space_15_lc_data(63 downto 32),
          mtag => memory_space_15_lc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_477_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_477_load_0_req_0;
      ptr_deref_477_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_477_load_0_req_1;
      ptr_deref_477_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_477_word_address_0;
      ptr_deref_477_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_16_lr_req(0),
          mack => memory_space_16_lr_ack(0),
          maddr => memory_space_16_lr_addr(0 downto 0),
          mtag => memory_space_16_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_16_lc_req(0),
          mack => memory_space_16_lc_ack(0),
          mdata => memory_space_16_lc_data(31 downto 0),
          mtag => memory_space_16_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_494_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_494_load_0_req_0;
      ptr_deref_494_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_494_load_0_req_1;
      ptr_deref_494_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_494_word_address_0;
      ptr_deref_494_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_15_lr_req(0),
          mack => memory_space_15_lr_ack(0),
          maddr => memory_space_15_lr_addr(0 downto 0),
          mtag => memory_space_15_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_15_lc_req(0),
          mack => memory_space_15_lc_ack(0),
          mdata => memory_space_15_lc_data(31 downto 0),
          mtag => memory_space_15_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : ptr_deref_441_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_441_store_0_req_0;
      ptr_deref_441_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_441_store_0_req_1;
      ptr_deref_441_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_441_word_address_0;
      data_in <= ptr_deref_441_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_15_sr_req(0),
          mack => memory_space_15_sr_ack(0),
          maddr => memory_space_15_sr_addr(0 downto 0),
          mdata => memory_space_15_sr_data(31 downto 0),
          mtag => memory_space_15_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_15_sc_req(0),
          mack => memory_space_15_sc_ack(0),
          mtag => memory_space_15_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_472_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_472_store_0_req_0;
      ptr_deref_472_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_472_store_0_req_1;
      ptr_deref_472_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_472_word_address_0;
      data_in <= ptr_deref_472_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_16_sr_req(0),
          mack => memory_space_16_sr_ack(0),
          maddr => memory_space_16_sr_addr(0 downto 0),
          mdata => memory_space_16_sr_data(31 downto 0),
          mtag => memory_space_16_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_16_sc_req(0),
          mack => memory_space_16_sc_ack(0),
          mtag => memory_space_16_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_489_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_489_store_0_req_0;
      ptr_deref_489_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_489_store_0_req_1;
      ptr_deref_489_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_489_word_address_0;
      data_in <= ptr_deref_489_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(2 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : simple_obj_ref_433_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_433_inst_req_0;
      simple_obj_ref_433_inst_ack_0 <= ack(0);
      simple_obj_ref_433_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_get_pipe_read_req(0),
          oack => free_queue_get_pipe_read_ack(0),
          odata => free_queue_get_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_468_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_468_inst_req_0;
      simple_obj_ref_468_inst_ack_0 <= ack(0);
      simple_obj_ref_468_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => input_data_pipe_read_req(0),
          oack => input_data_pipe_read_ack(0),
          odata => input_data_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_423_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_423_inst_req_0;
      simple_obj_ref_423_inst_ack_0 <= ack(0);
      data_in <= type_cast_425_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_505_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_505_inst_req_0;
      simple_obj_ref_505_inst_ack_0 <= ack(0);
      data_in <= type_cast_507_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => foo_in_pipe_write_req(0),
          oack => foo_in_pipe_write_ack(0),
          odata => foo_in_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  RegisterBank_memory_space_15: register_bank -- 
    generic map(-- 
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_15_lr_addr,
      lr_req_in => memory_space_15_lr_req,
      lr_ack_out => memory_space_15_lr_ack,
      lr_tag_in => memory_space_15_lr_tag,
      lc_req_in => memory_space_15_lc_req,
      lc_ack_out => memory_space_15_lc_ack,
      lc_data_out => memory_space_15_lc_data,
      lc_tag_out => memory_space_15_lc_tag,
      sr_addr_in => memory_space_15_sr_addr,
      sr_data_in => memory_space_15_sr_data,
      sr_req_in => memory_space_15_sr_req,
      sr_ack_out => memory_space_15_sr_ack,
      sr_tag_in => memory_space_15_sr_tag,
      sc_req_in=> memory_space_15_sc_req,
      sc_ack_out => memory_space_15_sc_ack,
      sc_tag_out => memory_space_15_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_16: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_16_lr_addr,
      lr_req_in => memory_space_16_lr_req,
      lr_ack_out => memory_space_16_lr_ack,
      lr_tag_in => memory_space_16_lr_tag,
      lc_req_in => memory_space_16_lc_req,
      lc_ack_out => memory_space_16_lc_ack,
      lc_data_out => memory_space_16_lc_data,
      lc_tag_out => memory_space_16_lc_tag,
      sr_addr_in => memory_space_16_sr_addr,
      sr_data_in => memory_space_16_sr_data,
      sr_req_in => memory_space_16_sr_req,
      sr_ack_out => memory_space_16_sr_ack,
      sr_tag_in => memory_space_16_sr_tag,
      sc_req_in=> memory_space_16_sc_req,
      sc_ack_out => memory_space_16_sc_ack,
      sc_tag_out => memory_space_16_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity mem_load_x_x is -- 
  port ( -- 
    address : in  std_logic_vector(31 downto 0);
    data : out  std_logic_vector(7 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity mem_load_x_x;
architecture Default of mem_load_x_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_13_load_0_ack_0 : boolean;
  signal binary_12_inst_req_0 : boolean;
  signal array_obj_ref_13_gather_scatter_ack_0 : boolean;
  signal binary_10_inst_ack_1 : boolean;
  signal array_obj_ref_13_load_0_req_0 : boolean;
  signal array_obj_ref_13_load_0_req_1 : boolean;
  signal binary_10_inst_req_1 : boolean;
  signal array_obj_ref_13_offset_inst_req_0 : boolean;
  signal array_obj_ref_13_offset_inst_ack_0 : boolean;
  signal array_obj_ref_13_gather_scatter_req_0 : boolean;
  signal binary_10_inst_ack_0 : boolean;
  signal binary_10_inst_req_0 : boolean;
  signal array_obj_ref_13_index_0_rename_req_0 : boolean;
  signal array_obj_ref_13_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_13_load_0_ack_1 : boolean;
  signal array_obj_ref_13_index_0_rename_ack_0 : boolean;
  signal binary_12_inst_ack_0 : boolean;
  signal binary_12_inst_req_1 : boolean;
  signal array_obj_ref_13_root_address_inst_req_0 : boolean;
  signal binary_12_inst_ack_1 : boolean;
  signal array_obj_ref_13_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_13_addr_0_req_0 : boolean;
  signal array_obj_ref_13_addr_0_ack_0 : boolean;
  signal array_obj_ref_13_index_0_resize_req_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  mem_load_x_xx_xCP_2275: Block -- control-path 
    signal mem_load_x_xx_xCP_2275_start: Boolean;
    signal Xentry_2276_symbol: Boolean;
    signal Xexit_2277_symbol: Boolean;
    signal assign_stmt_14_2278_symbol : Boolean;
    -- 
  begin -- 
    mem_load_x_xx_xCP_2275_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_2276_symbol  <= mem_load_x_xx_xCP_2275_start; -- transition $entry
    assign_stmt_14_2278: Block -- assign_stmt_14 
      signal assign_stmt_14_2278_start: Boolean;
      signal Xentry_2279_symbol: Boolean;
      signal Xexit_2280_symbol: Boolean;
      signal assign_stmt_14_active_x_x2281_symbol : Boolean;
      signal assign_stmt_14_completed_x_x2282_symbol : Boolean;
      signal array_obj_ref_13_trigger_x_x2283_symbol : Boolean;
      signal array_obj_ref_13_active_x_x2284_symbol : Boolean;
      signal array_obj_ref_13_root_address_calculated_2285_symbol : Boolean;
      signal array_obj_ref_13_word_address_calculated_2286_symbol : Boolean;
      signal array_obj_ref_13_indices_scaled_2287_symbol : Boolean;
      signal array_obj_ref_13_offset_calculated_2288_symbol : Boolean;
      signal array_obj_ref_13_index_computed_0_2289_symbol : Boolean;
      signal array_obj_ref_13_index_resized_0_2290_symbol : Boolean;
      signal binary_12_active_x_x2291_symbol : Boolean;
      signal binary_12_trigger_x_x2292_symbol : Boolean;
      signal binary_10_active_x_x2293_symbol : Boolean;
      signal binary_10_trigger_x_x2294_symbol : Boolean;
      signal simple_obj_ref_8_complete_2295_symbol : Boolean;
      signal binary_10_complete_2296_symbol : Boolean;
      signal binary_12_complete_2303_symbol : Boolean;
      signal array_obj_ref_13_index_resize_0_2310_symbol : Boolean;
      signal array_obj_ref_13_index_scale_0_2315_symbol : Boolean;
      signal array_obj_ref_13_add_indices_2320_symbol : Boolean;
      signal array_obj_ref_13_base_plus_offset_2325_symbol : Boolean;
      signal array_obj_ref_13_word_addrgen_2330_symbol : Boolean;
      signal array_obj_ref_13_request_2335_symbol : Boolean;
      signal array_obj_ref_13_complete_2346_symbol : Boolean;
      -- 
    begin -- 
      assign_stmt_14_2278_start <= Xentry_2276_symbol; -- control passed to block
      Xentry_2279_symbol  <= assign_stmt_14_2278_start; -- transition assign_stmt_14/$entry
      assign_stmt_14_active_x_x2281_symbol <= array_obj_ref_13_complete_2346_symbol; -- transition assign_stmt_14/assign_stmt_14_active_
      assign_stmt_14_completed_x_x2282_symbol <= assign_stmt_14_active_x_x2281_symbol; -- transition assign_stmt_14/assign_stmt_14_completed_
      array_obj_ref_13_trigger_x_x2283_symbol <= array_obj_ref_13_word_address_calculated_2286_symbol; -- transition assign_stmt_14/array_obj_ref_13_trigger_
      array_obj_ref_13_active_x_x2284_symbol <= array_obj_ref_13_request_2335_symbol; -- transition assign_stmt_14/array_obj_ref_13_active_
      array_obj_ref_13_root_address_calculated_2285_symbol <= array_obj_ref_13_base_plus_offset_2325_symbol; -- transition assign_stmt_14/array_obj_ref_13_root_address_calculated
      array_obj_ref_13_word_address_calculated_2286_symbol <= array_obj_ref_13_word_addrgen_2330_symbol; -- transition assign_stmt_14/array_obj_ref_13_word_address_calculated
      array_obj_ref_13_indices_scaled_2287_symbol <= array_obj_ref_13_index_scale_0_2315_symbol; -- transition assign_stmt_14/array_obj_ref_13_indices_scaled
      array_obj_ref_13_offset_calculated_2288_symbol <= array_obj_ref_13_add_indices_2320_symbol; -- transition assign_stmt_14/array_obj_ref_13_offset_calculated
      array_obj_ref_13_index_computed_0_2289_symbol <= binary_12_complete_2303_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_computed_0
      array_obj_ref_13_index_resized_0_2290_symbol <= array_obj_ref_13_index_resize_0_2310_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_resized_0
      binary_12_active_x_x2291_block : Block -- non-trivial join transition assign_stmt_14/binary_12_active_ 
        signal binary_12_active_x_x2291_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_12_active_x_x2291_predecessors(0) <= binary_12_trigger_x_x2292_symbol;
        binary_12_active_x_x2291_predecessors(1) <= binary_10_complete_2296_symbol;
        binary_12_active_x_x2291_join: join -- 
          port map( -- 
            preds => binary_12_active_x_x2291_predecessors,
            symbol_out => binary_12_active_x_x2291_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_14/binary_12_active_
      binary_12_trigger_x_x2292_symbol <= Xentry_2279_symbol; -- transition assign_stmt_14/binary_12_trigger_
      binary_10_active_x_x2293_block : Block -- non-trivial join transition assign_stmt_14/binary_10_active_ 
        signal binary_10_active_x_x2293_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_10_active_x_x2293_predecessors(0) <= binary_10_trigger_x_x2294_symbol;
        binary_10_active_x_x2293_predecessors(1) <= simple_obj_ref_8_complete_2295_symbol;
        binary_10_active_x_x2293_join: join -- 
          port map( -- 
            preds => binary_10_active_x_x2293_predecessors,
            symbol_out => binary_10_active_x_x2293_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_14/binary_10_active_
      binary_10_trigger_x_x2294_symbol <= Xentry_2279_symbol; -- transition assign_stmt_14/binary_10_trigger_
      simple_obj_ref_8_complete_2295_symbol <= Xentry_2279_symbol; -- transition assign_stmt_14/simple_obj_ref_8_complete
      binary_10_complete_2296: Block -- assign_stmt_14/binary_10_complete 
        signal binary_10_complete_2296_start: Boolean;
        signal Xentry_2297_symbol: Boolean;
        signal Xexit_2298_symbol: Boolean;
        signal rr_2299_symbol : Boolean;
        signal ra_2300_symbol : Boolean;
        signal cr_2301_symbol : Boolean;
        signal ca_2302_symbol : Boolean;
        -- 
      begin -- 
        binary_10_complete_2296_start <= binary_10_active_x_x2293_symbol; -- control passed to block
        Xentry_2297_symbol  <= binary_10_complete_2296_start; -- transition assign_stmt_14/binary_10_complete/$entry
        rr_2299_symbol <= Xentry_2297_symbol; -- transition assign_stmt_14/binary_10_complete/rr
        binary_10_inst_req_0 <= rr_2299_symbol; -- link to DP
        ra_2300_symbol <= binary_10_inst_ack_0; -- transition assign_stmt_14/binary_10_complete/ra
        cr_2301_symbol <= ra_2300_symbol; -- transition assign_stmt_14/binary_10_complete/cr
        binary_10_inst_req_1 <= cr_2301_symbol; -- link to DP
        ca_2302_symbol <= binary_10_inst_ack_1; -- transition assign_stmt_14/binary_10_complete/ca
        Xexit_2298_symbol <= ca_2302_symbol; -- transition assign_stmt_14/binary_10_complete/$exit
        binary_10_complete_2296_symbol <= Xexit_2298_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/binary_10_complete
      binary_12_complete_2303: Block -- assign_stmt_14/binary_12_complete 
        signal binary_12_complete_2303_start: Boolean;
        signal Xentry_2304_symbol: Boolean;
        signal Xexit_2305_symbol: Boolean;
        signal rr_2306_symbol : Boolean;
        signal ra_2307_symbol : Boolean;
        signal cr_2308_symbol : Boolean;
        signal ca_2309_symbol : Boolean;
        -- 
      begin -- 
        binary_12_complete_2303_start <= binary_12_active_x_x2291_symbol; -- control passed to block
        Xentry_2304_symbol  <= binary_12_complete_2303_start; -- transition assign_stmt_14/binary_12_complete/$entry
        rr_2306_symbol <= Xentry_2304_symbol; -- transition assign_stmt_14/binary_12_complete/rr
        binary_12_inst_req_0 <= rr_2306_symbol; -- link to DP
        ra_2307_symbol <= binary_12_inst_ack_0; -- transition assign_stmt_14/binary_12_complete/ra
        cr_2308_symbol <= ra_2307_symbol; -- transition assign_stmt_14/binary_12_complete/cr
        binary_12_inst_req_1 <= cr_2308_symbol; -- link to DP
        ca_2309_symbol <= binary_12_inst_ack_1; -- transition assign_stmt_14/binary_12_complete/ca
        Xexit_2305_symbol <= ca_2309_symbol; -- transition assign_stmt_14/binary_12_complete/$exit
        binary_12_complete_2303_symbol <= Xexit_2305_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/binary_12_complete
      array_obj_ref_13_index_resize_0_2310: Block -- assign_stmt_14/array_obj_ref_13_index_resize_0 
        signal array_obj_ref_13_index_resize_0_2310_start: Boolean;
        signal Xentry_2311_symbol: Boolean;
        signal Xexit_2312_symbol: Boolean;
        signal index_resize_req_2313_symbol : Boolean;
        signal index_resize_ack_2314_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_index_resize_0_2310_start <= array_obj_ref_13_index_computed_0_2289_symbol; -- control passed to block
        Xentry_2311_symbol  <= array_obj_ref_13_index_resize_0_2310_start; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/$entry
        index_resize_req_2313_symbol <= Xentry_2311_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/index_resize_req
        array_obj_ref_13_index_0_resize_req_0 <= index_resize_req_2313_symbol; -- link to DP
        index_resize_ack_2314_symbol <= array_obj_ref_13_index_0_resize_ack_0; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/index_resize_ack
        Xexit_2312_symbol <= index_resize_ack_2314_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_resize_0/$exit
        array_obj_ref_13_index_resize_0_2310_symbol <= Xexit_2312_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_index_resize_0
      array_obj_ref_13_index_scale_0_2315: Block -- assign_stmt_14/array_obj_ref_13_index_scale_0 
        signal array_obj_ref_13_index_scale_0_2315_start: Boolean;
        signal Xentry_2316_symbol: Boolean;
        signal Xexit_2317_symbol: Boolean;
        signal scale_rename_req_2318_symbol : Boolean;
        signal scale_rename_ack_2319_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_index_scale_0_2315_start <= array_obj_ref_13_index_resized_0_2290_symbol; -- control passed to block
        Xentry_2316_symbol  <= array_obj_ref_13_index_scale_0_2315_start; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/$entry
        scale_rename_req_2318_symbol <= Xentry_2316_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/scale_rename_req
        array_obj_ref_13_index_0_rename_req_0 <= scale_rename_req_2318_symbol; -- link to DP
        scale_rename_ack_2319_symbol <= array_obj_ref_13_index_0_rename_ack_0; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/scale_rename_ack
        Xexit_2317_symbol <= scale_rename_ack_2319_symbol; -- transition assign_stmt_14/array_obj_ref_13_index_scale_0/$exit
        array_obj_ref_13_index_scale_0_2315_symbol <= Xexit_2317_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_index_scale_0
      array_obj_ref_13_add_indices_2320: Block -- assign_stmt_14/array_obj_ref_13_add_indices 
        signal array_obj_ref_13_add_indices_2320_start: Boolean;
        signal Xentry_2321_symbol: Boolean;
        signal Xexit_2322_symbol: Boolean;
        signal final_index_req_2323_symbol : Boolean;
        signal final_index_ack_2324_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_add_indices_2320_start <= array_obj_ref_13_indices_scaled_2287_symbol; -- control passed to block
        Xentry_2321_symbol  <= array_obj_ref_13_add_indices_2320_start; -- transition assign_stmt_14/array_obj_ref_13_add_indices/$entry
        final_index_req_2323_symbol <= Xentry_2321_symbol; -- transition assign_stmt_14/array_obj_ref_13_add_indices/final_index_req
        array_obj_ref_13_offset_inst_req_0 <= final_index_req_2323_symbol; -- link to DP
        final_index_ack_2324_symbol <= array_obj_ref_13_offset_inst_ack_0; -- transition assign_stmt_14/array_obj_ref_13_add_indices/final_index_ack
        Xexit_2322_symbol <= final_index_ack_2324_symbol; -- transition assign_stmt_14/array_obj_ref_13_add_indices/$exit
        array_obj_ref_13_add_indices_2320_symbol <= Xexit_2322_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_add_indices
      array_obj_ref_13_base_plus_offset_2325: Block -- assign_stmt_14/array_obj_ref_13_base_plus_offset 
        signal array_obj_ref_13_base_plus_offset_2325_start: Boolean;
        signal Xentry_2326_symbol: Boolean;
        signal Xexit_2327_symbol: Boolean;
        signal sum_rename_req_2328_symbol : Boolean;
        signal sum_rename_ack_2329_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_base_plus_offset_2325_start <= array_obj_ref_13_offset_calculated_2288_symbol; -- control passed to block
        Xentry_2326_symbol  <= array_obj_ref_13_base_plus_offset_2325_start; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/$entry
        sum_rename_req_2328_symbol <= Xentry_2326_symbol; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/sum_rename_req
        array_obj_ref_13_root_address_inst_req_0 <= sum_rename_req_2328_symbol; -- link to DP
        sum_rename_ack_2329_symbol <= array_obj_ref_13_root_address_inst_ack_0; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/sum_rename_ack
        Xexit_2327_symbol <= sum_rename_ack_2329_symbol; -- transition assign_stmt_14/array_obj_ref_13_base_plus_offset/$exit
        array_obj_ref_13_base_plus_offset_2325_symbol <= Xexit_2327_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_base_plus_offset
      array_obj_ref_13_word_addrgen_2330: Block -- assign_stmt_14/array_obj_ref_13_word_addrgen 
        signal array_obj_ref_13_word_addrgen_2330_start: Boolean;
        signal Xentry_2331_symbol: Boolean;
        signal Xexit_2332_symbol: Boolean;
        signal root_rename_req_2333_symbol : Boolean;
        signal root_rename_ack_2334_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_word_addrgen_2330_start <= array_obj_ref_13_root_address_calculated_2285_symbol; -- control passed to block
        Xentry_2331_symbol  <= array_obj_ref_13_word_addrgen_2330_start; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/$entry
        root_rename_req_2333_symbol <= Xentry_2331_symbol; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/root_rename_req
        array_obj_ref_13_addr_0_req_0 <= root_rename_req_2333_symbol; -- link to DP
        root_rename_ack_2334_symbol <= array_obj_ref_13_addr_0_ack_0; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/root_rename_ack
        Xexit_2332_symbol <= root_rename_ack_2334_symbol; -- transition assign_stmt_14/array_obj_ref_13_word_addrgen/$exit
        array_obj_ref_13_word_addrgen_2330_symbol <= Xexit_2332_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_word_addrgen
      array_obj_ref_13_request_2335: Block -- assign_stmt_14/array_obj_ref_13_request 
        signal array_obj_ref_13_request_2335_start: Boolean;
        signal Xentry_2336_symbol: Boolean;
        signal Xexit_2337_symbol: Boolean;
        signal word_access_2338_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_request_2335_start <= array_obj_ref_13_trigger_x_x2283_symbol; -- control passed to block
        Xentry_2336_symbol  <= array_obj_ref_13_request_2335_start; -- transition assign_stmt_14/array_obj_ref_13_request/$entry
        word_access_2338: Block -- assign_stmt_14/array_obj_ref_13_request/word_access 
          signal word_access_2338_start: Boolean;
          signal Xentry_2339_symbol: Boolean;
          signal Xexit_2340_symbol: Boolean;
          signal word_access_0_2341_symbol : Boolean;
          -- 
        begin -- 
          word_access_2338_start <= Xentry_2336_symbol; -- control passed to block
          Xentry_2339_symbol  <= word_access_2338_start; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/$entry
          word_access_0_2341: Block -- assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0 
            signal word_access_0_2341_start: Boolean;
            signal Xentry_2342_symbol: Boolean;
            signal Xexit_2343_symbol: Boolean;
            signal rr_2344_symbol : Boolean;
            signal ra_2345_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_2341_start <= Xentry_2339_symbol; -- control passed to block
            Xentry_2342_symbol  <= word_access_0_2341_start; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/$entry
            rr_2344_symbol <= Xentry_2342_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/rr
            array_obj_ref_13_load_0_req_0 <= rr_2344_symbol; -- link to DP
            ra_2345_symbol <= array_obj_ref_13_load_0_ack_0; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/ra
            Xexit_2343_symbol <= ra_2345_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0/$exit
            word_access_0_2341_symbol <= Xexit_2343_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_14/array_obj_ref_13_request/word_access/word_access_0
          Xexit_2340_symbol <= word_access_0_2341_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/word_access/$exit
          word_access_2338_symbol <= Xexit_2340_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_14/array_obj_ref_13_request/word_access
        Xexit_2337_symbol <= word_access_2338_symbol; -- transition assign_stmt_14/array_obj_ref_13_request/$exit
        array_obj_ref_13_request_2335_symbol <= Xexit_2337_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_request
      array_obj_ref_13_complete_2346: Block -- assign_stmt_14/array_obj_ref_13_complete 
        signal array_obj_ref_13_complete_2346_start: Boolean;
        signal Xentry_2347_symbol: Boolean;
        signal Xexit_2348_symbol: Boolean;
        signal word_access_2349_symbol : Boolean;
        signal merge_req_2357_symbol : Boolean;
        signal merge_ack_2358_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_13_complete_2346_start <= array_obj_ref_13_active_x_x2284_symbol; -- control passed to block
        Xentry_2347_symbol  <= array_obj_ref_13_complete_2346_start; -- transition assign_stmt_14/array_obj_ref_13_complete/$entry
        word_access_2349: Block -- assign_stmt_14/array_obj_ref_13_complete/word_access 
          signal word_access_2349_start: Boolean;
          signal Xentry_2350_symbol: Boolean;
          signal Xexit_2351_symbol: Boolean;
          signal word_access_0_2352_symbol : Boolean;
          -- 
        begin -- 
          word_access_2349_start <= Xentry_2347_symbol; -- control passed to block
          Xentry_2350_symbol  <= word_access_2349_start; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/$entry
          word_access_0_2352: Block -- assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0 
            signal word_access_0_2352_start: Boolean;
            signal Xentry_2353_symbol: Boolean;
            signal Xexit_2354_symbol: Boolean;
            signal cr_2355_symbol : Boolean;
            signal ca_2356_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_2352_start <= Xentry_2350_symbol; -- control passed to block
            Xentry_2353_symbol  <= word_access_0_2352_start; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/$entry
            cr_2355_symbol <= Xentry_2353_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/cr
            array_obj_ref_13_load_0_req_1 <= cr_2355_symbol; -- link to DP
            ca_2356_symbol <= array_obj_ref_13_load_0_ack_1; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/ca
            Xexit_2354_symbol <= ca_2356_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0/$exit
            word_access_0_2352_symbol <= Xexit_2354_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_14/array_obj_ref_13_complete/word_access/word_access_0
          Xexit_2351_symbol <= word_access_0_2352_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/word_access/$exit
          word_access_2349_symbol <= Xexit_2351_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_14/array_obj_ref_13_complete/word_access
        merge_req_2357_symbol <= word_access_2349_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/merge_req
        array_obj_ref_13_gather_scatter_req_0 <= merge_req_2357_symbol; -- link to DP
        merge_ack_2358_symbol <= array_obj_ref_13_gather_scatter_ack_0; -- transition assign_stmt_14/array_obj_ref_13_complete/merge_ack
        Xexit_2348_symbol <= merge_ack_2358_symbol; -- transition assign_stmt_14/array_obj_ref_13_complete/$exit
        array_obj_ref_13_complete_2346_symbol <= Xexit_2348_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_14/array_obj_ref_13_complete
      Xexit_2280_symbol <= assign_stmt_14_completed_x_x2282_symbol; -- transition assign_stmt_14/$exit
      assign_stmt_14_2278_symbol <= Xexit_2280_symbol; -- control passed from block 
      -- 
    end Block; -- assign_stmt_14
    Xexit_2277_symbol <= assign_stmt_14_2278_symbol; -- transition $exit
    fin  <=  '1' when Xexit_2277_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_13_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_13_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_word_address_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_13_word_offset_0 : std_logic_vector(0 downto 0);
    signal binary_10_wire : std_logic_vector(31 downto 0);
    signal binary_12_resized : std_logic_vector(0 downto 0);
    signal binary_12_scaled : std_logic_vector(0 downto 0);
    signal binary_12_wire : std_logic_vector(31 downto 0);
    signal expr_11_wire_constant : std_logic_vector(31 downto 0);
    signal expr_9_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_13_offset_scale_factor_0 <= "1";
    array_obj_ref_13_resized_base_address <= "0";
    array_obj_ref_13_word_offset_0 <= "0";
    expr_11_wire_constant <= "00000000000000000000000000000000";
    expr_9_wire_constant <= "00000000000000000000000000000001";
    array_obj_ref_13_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 1) -- 
      port map( din => binary_12_wire, dout => binary_12_resized, req => array_obj_ref_13_index_0_resize_req_0, ack => array_obj_ref_13_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_13_offset_inst: RegisterBase generic map(in_data_width => 1,out_data_width => 1) -- 
      port map( din => binary_12_scaled, dout => array_obj_ref_13_final_offset, req => array_obj_ref_13_offset_inst_req_0, ack => array_obj_ref_13_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_13_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_13_addr_0_ack_0 <= array_obj_ref_13_addr_0_req_0;
      aggregated_sig <= array_obj_ref_13_root_address;
      array_obj_ref_13_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_13_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_13_gather_scatter_ack_0 <= array_obj_ref_13_gather_scatter_req_0;
      aggregated_sig <= array_obj_ref_13_data_0;
      data <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_13_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_13_index_0_rename_ack_0 <= array_obj_ref_13_index_0_rename_req_0;
      aggregated_sig <= binary_12_resized;
      binary_12_scaled <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_13_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_13_root_address_inst_ack_0 <= array_obj_ref_13_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_13_final_offset;
      array_obj_ref_13_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    -- shared split operator group (0) : binary_10_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= address;
      binary_10_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_10_inst_req_0,
          ackL => binary_10_inst_ack_0,
          reqR => binary_10_inst_req_1,
          ackR => binary_10_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_12_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_10_wire;
      binary_12_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_12_inst_req_0,
          ackL => binary_12_inst_ack_0,
          reqR => binary_12_inst_req_1,
          ackR => binary_12_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared load operator group (0) : array_obj_ref_13_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_13_load_0_req_0;
      array_obj_ref_13_load_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_13_load_0_req_1;
      array_obj_ref_13_load_0_ack_1 <= ackR(0);
      data_in <= array_obj_ref_13_word_address_0;
      array_obj_ref_13_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 1,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(7 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity mem_store_x_x is -- 
  port ( -- 
    address : in  std_logic_vector(31 downto 0);
    data : in  std_logic_vector(7 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity mem_store_x_x;
architecture Default of mem_store_x_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal binary_21_inst_req_0 : boolean;
  signal array_obj_ref_24_store_0_ack_1 : boolean;
  signal binary_21_inst_req_1 : boolean;
  signal array_obj_ref_24_store_0_req_1 : boolean;
  signal binary_23_inst_ack_1 : boolean;
  signal array_obj_ref_24_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_24_index_0_rename_req_0 : boolean;
  signal array_obj_ref_24_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_24_offset_inst_req_0 : boolean;
  signal array_obj_ref_24_offset_inst_ack_0 : boolean;
  signal array_obj_ref_24_store_0_ack_0 : boolean;
  signal array_obj_ref_24_addr_0_ack_0 : boolean;
  signal array_obj_ref_24_store_0_req_0 : boolean;
  signal array_obj_ref_24_index_0_rename_ack_0 : boolean;
  signal binary_23_inst_ack_0 : boolean;
  signal array_obj_ref_24_index_0_resize_req_0 : boolean;
  signal binary_23_inst_req_1 : boolean;
  signal array_obj_ref_24_addr_0_req_0 : boolean;
  signal array_obj_ref_24_root_address_inst_req_0 : boolean;
  signal array_obj_ref_24_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_24_gather_scatter_req_0 : boolean;
  signal binary_21_inst_ack_0 : boolean;
  signal binary_21_inst_ack_1 : boolean;
  signal binary_23_inst_req_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  mem_store_x_xx_xCP_2359: Block -- control-path 
    signal mem_store_x_xx_xCP_2359_start: Boolean;
    signal Xentry_2360_symbol: Boolean;
    signal Xexit_2361_symbol: Boolean;
    signal assign_stmt_26_2362_symbol : Boolean;
    -- 
  begin -- 
    mem_store_x_xx_xCP_2359_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_2360_symbol  <= mem_store_x_xx_xCP_2359_start; -- transition $entry
    assign_stmt_26_2362: Block -- assign_stmt_26 
      signal assign_stmt_26_2362_start: Boolean;
      signal Xentry_2363_symbol: Boolean;
      signal Xexit_2364_symbol: Boolean;
      signal assign_stmt_26_active_x_x2365_symbol : Boolean;
      signal assign_stmt_26_completed_x_x2366_symbol : Boolean;
      signal simple_obj_ref_25_complete_2367_symbol : Boolean;
      signal array_obj_ref_24_trigger_x_x2368_symbol : Boolean;
      signal array_obj_ref_24_active_x_x2369_symbol : Boolean;
      signal array_obj_ref_24_root_address_calculated_2370_symbol : Boolean;
      signal array_obj_ref_24_word_address_calculated_2371_symbol : Boolean;
      signal array_obj_ref_24_indices_scaled_2372_symbol : Boolean;
      signal array_obj_ref_24_offset_calculated_2373_symbol : Boolean;
      signal array_obj_ref_24_index_computed_0_2374_symbol : Boolean;
      signal array_obj_ref_24_index_resized_0_2375_symbol : Boolean;
      signal binary_23_active_x_x2376_symbol : Boolean;
      signal binary_23_trigger_x_x2377_symbol : Boolean;
      signal binary_21_active_x_x2378_symbol : Boolean;
      signal binary_21_trigger_x_x2379_symbol : Boolean;
      signal simple_obj_ref_19_complete_2380_symbol : Boolean;
      signal binary_21_complete_2381_symbol : Boolean;
      signal binary_23_complete_2388_symbol : Boolean;
      signal array_obj_ref_24_index_resize_0_2395_symbol : Boolean;
      signal array_obj_ref_24_index_scale_0_2400_symbol : Boolean;
      signal array_obj_ref_24_add_indices_2405_symbol : Boolean;
      signal array_obj_ref_24_base_plus_offset_2410_symbol : Boolean;
      signal array_obj_ref_24_word_addrgen_2415_symbol : Boolean;
      signal array_obj_ref_24_request_2420_symbol : Boolean;
      signal array_obj_ref_24_complete_2433_symbol : Boolean;
      -- 
    begin -- 
      assign_stmt_26_2362_start <= Xentry_2360_symbol; -- control passed to block
      Xentry_2363_symbol  <= assign_stmt_26_2362_start; -- transition assign_stmt_26/$entry
      assign_stmt_26_active_x_x2365_symbol <= simple_obj_ref_25_complete_2367_symbol; -- transition assign_stmt_26/assign_stmt_26_active_
      assign_stmt_26_completed_x_x2366_symbol <= array_obj_ref_24_complete_2433_symbol; -- transition assign_stmt_26/assign_stmt_26_completed_
      simple_obj_ref_25_complete_2367_symbol <= Xentry_2363_symbol; -- transition assign_stmt_26/simple_obj_ref_25_complete
      array_obj_ref_24_trigger_x_x2368_block : Block -- non-trivial join transition assign_stmt_26/array_obj_ref_24_trigger_ 
        signal array_obj_ref_24_trigger_x_x2368_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        array_obj_ref_24_trigger_x_x2368_predecessors(0) <= array_obj_ref_24_word_address_calculated_2371_symbol;
        array_obj_ref_24_trigger_x_x2368_predecessors(1) <= assign_stmt_26_active_x_x2365_symbol;
        array_obj_ref_24_trigger_x_x2368_join: join -- 
          port map( -- 
            preds => array_obj_ref_24_trigger_x_x2368_predecessors,
            symbol_out => array_obj_ref_24_trigger_x_x2368_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_26/array_obj_ref_24_trigger_
      array_obj_ref_24_active_x_x2369_symbol <= array_obj_ref_24_request_2420_symbol; -- transition assign_stmt_26/array_obj_ref_24_active_
      array_obj_ref_24_root_address_calculated_2370_symbol <= array_obj_ref_24_base_plus_offset_2410_symbol; -- transition assign_stmt_26/array_obj_ref_24_root_address_calculated
      array_obj_ref_24_word_address_calculated_2371_symbol <= array_obj_ref_24_word_addrgen_2415_symbol; -- transition assign_stmt_26/array_obj_ref_24_word_address_calculated
      array_obj_ref_24_indices_scaled_2372_symbol <= array_obj_ref_24_index_scale_0_2400_symbol; -- transition assign_stmt_26/array_obj_ref_24_indices_scaled
      array_obj_ref_24_offset_calculated_2373_symbol <= array_obj_ref_24_add_indices_2405_symbol; -- transition assign_stmt_26/array_obj_ref_24_offset_calculated
      array_obj_ref_24_index_computed_0_2374_symbol <= binary_23_complete_2388_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_computed_0
      array_obj_ref_24_index_resized_0_2375_symbol <= array_obj_ref_24_index_resize_0_2395_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_resized_0
      binary_23_active_x_x2376_block : Block -- non-trivial join transition assign_stmt_26/binary_23_active_ 
        signal binary_23_active_x_x2376_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_23_active_x_x2376_predecessors(0) <= binary_23_trigger_x_x2377_symbol;
        binary_23_active_x_x2376_predecessors(1) <= binary_21_complete_2381_symbol;
        binary_23_active_x_x2376_join: join -- 
          port map( -- 
            preds => binary_23_active_x_x2376_predecessors,
            symbol_out => binary_23_active_x_x2376_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_26/binary_23_active_
      binary_23_trigger_x_x2377_symbol <= Xentry_2363_symbol; -- transition assign_stmt_26/binary_23_trigger_
      binary_21_active_x_x2378_block : Block -- non-trivial join transition assign_stmt_26/binary_21_active_ 
        signal binary_21_active_x_x2378_predecessors: BooleanArray(1 downto 0);
        -- 
      begin -- 
        binary_21_active_x_x2378_predecessors(0) <= binary_21_trigger_x_x2379_symbol;
        binary_21_active_x_x2378_predecessors(1) <= simple_obj_ref_19_complete_2380_symbol;
        binary_21_active_x_x2378_join: join -- 
          port map( -- 
            preds => binary_21_active_x_x2378_predecessors,
            symbol_out => binary_21_active_x_x2378_symbol,
            clk => clk,
            reset => reset); -- 
        -- 
      end Block; -- non-trivial join transition assign_stmt_26/binary_21_active_
      binary_21_trigger_x_x2379_symbol <= Xentry_2363_symbol; -- transition assign_stmt_26/binary_21_trigger_
      simple_obj_ref_19_complete_2380_symbol <= Xentry_2363_symbol; -- transition assign_stmt_26/simple_obj_ref_19_complete
      binary_21_complete_2381: Block -- assign_stmt_26/binary_21_complete 
        signal binary_21_complete_2381_start: Boolean;
        signal Xentry_2382_symbol: Boolean;
        signal Xexit_2383_symbol: Boolean;
        signal rr_2384_symbol : Boolean;
        signal ra_2385_symbol : Boolean;
        signal cr_2386_symbol : Boolean;
        signal ca_2387_symbol : Boolean;
        -- 
      begin -- 
        binary_21_complete_2381_start <= binary_21_active_x_x2378_symbol; -- control passed to block
        Xentry_2382_symbol  <= binary_21_complete_2381_start; -- transition assign_stmt_26/binary_21_complete/$entry
        rr_2384_symbol <= Xentry_2382_symbol; -- transition assign_stmt_26/binary_21_complete/rr
        binary_21_inst_req_0 <= rr_2384_symbol; -- link to DP
        ra_2385_symbol <= binary_21_inst_ack_0; -- transition assign_stmt_26/binary_21_complete/ra
        cr_2386_symbol <= ra_2385_symbol; -- transition assign_stmt_26/binary_21_complete/cr
        binary_21_inst_req_1 <= cr_2386_symbol; -- link to DP
        ca_2387_symbol <= binary_21_inst_ack_1; -- transition assign_stmt_26/binary_21_complete/ca
        Xexit_2383_symbol <= ca_2387_symbol; -- transition assign_stmt_26/binary_21_complete/$exit
        binary_21_complete_2381_symbol <= Xexit_2383_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/binary_21_complete
      binary_23_complete_2388: Block -- assign_stmt_26/binary_23_complete 
        signal binary_23_complete_2388_start: Boolean;
        signal Xentry_2389_symbol: Boolean;
        signal Xexit_2390_symbol: Boolean;
        signal rr_2391_symbol : Boolean;
        signal ra_2392_symbol : Boolean;
        signal cr_2393_symbol : Boolean;
        signal ca_2394_symbol : Boolean;
        -- 
      begin -- 
        binary_23_complete_2388_start <= binary_23_active_x_x2376_symbol; -- control passed to block
        Xentry_2389_symbol  <= binary_23_complete_2388_start; -- transition assign_stmt_26/binary_23_complete/$entry
        rr_2391_symbol <= Xentry_2389_symbol; -- transition assign_stmt_26/binary_23_complete/rr
        binary_23_inst_req_0 <= rr_2391_symbol; -- link to DP
        ra_2392_symbol <= binary_23_inst_ack_0; -- transition assign_stmt_26/binary_23_complete/ra
        cr_2393_symbol <= ra_2392_symbol; -- transition assign_stmt_26/binary_23_complete/cr
        binary_23_inst_req_1 <= cr_2393_symbol; -- link to DP
        ca_2394_symbol <= binary_23_inst_ack_1; -- transition assign_stmt_26/binary_23_complete/ca
        Xexit_2390_symbol <= ca_2394_symbol; -- transition assign_stmt_26/binary_23_complete/$exit
        binary_23_complete_2388_symbol <= Xexit_2390_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/binary_23_complete
      array_obj_ref_24_index_resize_0_2395: Block -- assign_stmt_26/array_obj_ref_24_index_resize_0 
        signal array_obj_ref_24_index_resize_0_2395_start: Boolean;
        signal Xentry_2396_symbol: Boolean;
        signal Xexit_2397_symbol: Boolean;
        signal index_resize_req_2398_symbol : Boolean;
        signal index_resize_ack_2399_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_index_resize_0_2395_start <= array_obj_ref_24_index_computed_0_2374_symbol; -- control passed to block
        Xentry_2396_symbol  <= array_obj_ref_24_index_resize_0_2395_start; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/$entry
        index_resize_req_2398_symbol <= Xentry_2396_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/index_resize_req
        array_obj_ref_24_index_0_resize_req_0 <= index_resize_req_2398_symbol; -- link to DP
        index_resize_ack_2399_symbol <= array_obj_ref_24_index_0_resize_ack_0; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/index_resize_ack
        Xexit_2397_symbol <= index_resize_ack_2399_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_resize_0/$exit
        array_obj_ref_24_index_resize_0_2395_symbol <= Xexit_2397_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_index_resize_0
      array_obj_ref_24_index_scale_0_2400: Block -- assign_stmt_26/array_obj_ref_24_index_scale_0 
        signal array_obj_ref_24_index_scale_0_2400_start: Boolean;
        signal Xentry_2401_symbol: Boolean;
        signal Xexit_2402_symbol: Boolean;
        signal scale_rename_req_2403_symbol : Boolean;
        signal scale_rename_ack_2404_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_index_scale_0_2400_start <= array_obj_ref_24_index_resized_0_2375_symbol; -- control passed to block
        Xentry_2401_symbol  <= array_obj_ref_24_index_scale_0_2400_start; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/$entry
        scale_rename_req_2403_symbol <= Xentry_2401_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/scale_rename_req
        array_obj_ref_24_index_0_rename_req_0 <= scale_rename_req_2403_symbol; -- link to DP
        scale_rename_ack_2404_symbol <= array_obj_ref_24_index_0_rename_ack_0; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/scale_rename_ack
        Xexit_2402_symbol <= scale_rename_ack_2404_symbol; -- transition assign_stmt_26/array_obj_ref_24_index_scale_0/$exit
        array_obj_ref_24_index_scale_0_2400_symbol <= Xexit_2402_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_index_scale_0
      array_obj_ref_24_add_indices_2405: Block -- assign_stmt_26/array_obj_ref_24_add_indices 
        signal array_obj_ref_24_add_indices_2405_start: Boolean;
        signal Xentry_2406_symbol: Boolean;
        signal Xexit_2407_symbol: Boolean;
        signal final_index_req_2408_symbol : Boolean;
        signal final_index_ack_2409_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_add_indices_2405_start <= array_obj_ref_24_indices_scaled_2372_symbol; -- control passed to block
        Xentry_2406_symbol  <= array_obj_ref_24_add_indices_2405_start; -- transition assign_stmt_26/array_obj_ref_24_add_indices/$entry
        final_index_req_2408_symbol <= Xentry_2406_symbol; -- transition assign_stmt_26/array_obj_ref_24_add_indices/final_index_req
        array_obj_ref_24_offset_inst_req_0 <= final_index_req_2408_symbol; -- link to DP
        final_index_ack_2409_symbol <= array_obj_ref_24_offset_inst_ack_0; -- transition assign_stmt_26/array_obj_ref_24_add_indices/final_index_ack
        Xexit_2407_symbol <= final_index_ack_2409_symbol; -- transition assign_stmt_26/array_obj_ref_24_add_indices/$exit
        array_obj_ref_24_add_indices_2405_symbol <= Xexit_2407_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_add_indices
      array_obj_ref_24_base_plus_offset_2410: Block -- assign_stmt_26/array_obj_ref_24_base_plus_offset 
        signal array_obj_ref_24_base_plus_offset_2410_start: Boolean;
        signal Xentry_2411_symbol: Boolean;
        signal Xexit_2412_symbol: Boolean;
        signal sum_rename_req_2413_symbol : Boolean;
        signal sum_rename_ack_2414_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_base_plus_offset_2410_start <= array_obj_ref_24_offset_calculated_2373_symbol; -- control passed to block
        Xentry_2411_symbol  <= array_obj_ref_24_base_plus_offset_2410_start; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/$entry
        sum_rename_req_2413_symbol <= Xentry_2411_symbol; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/sum_rename_req
        array_obj_ref_24_root_address_inst_req_0 <= sum_rename_req_2413_symbol; -- link to DP
        sum_rename_ack_2414_symbol <= array_obj_ref_24_root_address_inst_ack_0; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/sum_rename_ack
        Xexit_2412_symbol <= sum_rename_ack_2414_symbol; -- transition assign_stmt_26/array_obj_ref_24_base_plus_offset/$exit
        array_obj_ref_24_base_plus_offset_2410_symbol <= Xexit_2412_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_base_plus_offset
      array_obj_ref_24_word_addrgen_2415: Block -- assign_stmt_26/array_obj_ref_24_word_addrgen 
        signal array_obj_ref_24_word_addrgen_2415_start: Boolean;
        signal Xentry_2416_symbol: Boolean;
        signal Xexit_2417_symbol: Boolean;
        signal root_rename_req_2418_symbol : Boolean;
        signal root_rename_ack_2419_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_word_addrgen_2415_start <= array_obj_ref_24_root_address_calculated_2370_symbol; -- control passed to block
        Xentry_2416_symbol  <= array_obj_ref_24_word_addrgen_2415_start; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/$entry
        root_rename_req_2418_symbol <= Xentry_2416_symbol; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/root_rename_req
        array_obj_ref_24_addr_0_req_0 <= root_rename_req_2418_symbol; -- link to DP
        root_rename_ack_2419_symbol <= array_obj_ref_24_addr_0_ack_0; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/root_rename_ack
        Xexit_2417_symbol <= root_rename_ack_2419_symbol; -- transition assign_stmt_26/array_obj_ref_24_word_addrgen/$exit
        array_obj_ref_24_word_addrgen_2415_symbol <= Xexit_2417_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_word_addrgen
      array_obj_ref_24_request_2420: Block -- assign_stmt_26/array_obj_ref_24_request 
        signal array_obj_ref_24_request_2420_start: Boolean;
        signal Xentry_2421_symbol: Boolean;
        signal Xexit_2422_symbol: Boolean;
        signal split_req_2423_symbol : Boolean;
        signal split_ack_2424_symbol : Boolean;
        signal word_access_2425_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_request_2420_start <= array_obj_ref_24_trigger_x_x2368_symbol; -- control passed to block
        Xentry_2421_symbol  <= array_obj_ref_24_request_2420_start; -- transition assign_stmt_26/array_obj_ref_24_request/$entry
        split_req_2423_symbol <= Xentry_2421_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/split_req
        array_obj_ref_24_gather_scatter_req_0 <= split_req_2423_symbol; -- link to DP
        split_ack_2424_symbol <= array_obj_ref_24_gather_scatter_ack_0; -- transition assign_stmt_26/array_obj_ref_24_request/split_ack
        word_access_2425: Block -- assign_stmt_26/array_obj_ref_24_request/word_access 
          signal word_access_2425_start: Boolean;
          signal Xentry_2426_symbol: Boolean;
          signal Xexit_2427_symbol: Boolean;
          signal word_access_0_2428_symbol : Boolean;
          -- 
        begin -- 
          word_access_2425_start <= split_ack_2424_symbol; -- control passed to block
          Xentry_2426_symbol  <= word_access_2425_start; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/$entry
          word_access_0_2428: Block -- assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0 
            signal word_access_0_2428_start: Boolean;
            signal Xentry_2429_symbol: Boolean;
            signal Xexit_2430_symbol: Boolean;
            signal rr_2431_symbol : Boolean;
            signal ra_2432_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_2428_start <= Xentry_2426_symbol; -- control passed to block
            Xentry_2429_symbol  <= word_access_0_2428_start; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/$entry
            rr_2431_symbol <= Xentry_2429_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/rr
            array_obj_ref_24_store_0_req_0 <= rr_2431_symbol; -- link to DP
            ra_2432_symbol <= array_obj_ref_24_store_0_ack_0; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/ra
            Xexit_2430_symbol <= ra_2432_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0/$exit
            word_access_0_2428_symbol <= Xexit_2430_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_26/array_obj_ref_24_request/word_access/word_access_0
          Xexit_2427_symbol <= word_access_0_2428_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/word_access/$exit
          word_access_2425_symbol <= Xexit_2427_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_26/array_obj_ref_24_request/word_access
        Xexit_2422_symbol <= word_access_2425_symbol; -- transition assign_stmt_26/array_obj_ref_24_request/$exit
        array_obj_ref_24_request_2420_symbol <= Xexit_2422_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_request
      array_obj_ref_24_complete_2433: Block -- assign_stmt_26/array_obj_ref_24_complete 
        signal array_obj_ref_24_complete_2433_start: Boolean;
        signal Xentry_2434_symbol: Boolean;
        signal Xexit_2435_symbol: Boolean;
        signal word_access_2436_symbol : Boolean;
        -- 
      begin -- 
        array_obj_ref_24_complete_2433_start <= array_obj_ref_24_active_x_x2369_symbol; -- control passed to block
        Xentry_2434_symbol  <= array_obj_ref_24_complete_2433_start; -- transition assign_stmt_26/array_obj_ref_24_complete/$entry
        word_access_2436: Block -- assign_stmt_26/array_obj_ref_24_complete/word_access 
          signal word_access_2436_start: Boolean;
          signal Xentry_2437_symbol: Boolean;
          signal Xexit_2438_symbol: Boolean;
          signal word_access_0_2439_symbol : Boolean;
          -- 
        begin -- 
          word_access_2436_start <= Xentry_2434_symbol; -- control passed to block
          Xentry_2437_symbol  <= word_access_2436_start; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/$entry
          word_access_0_2439: Block -- assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0 
            signal word_access_0_2439_start: Boolean;
            signal Xentry_2440_symbol: Boolean;
            signal Xexit_2441_symbol: Boolean;
            signal cr_2442_symbol : Boolean;
            signal ca_2443_symbol : Boolean;
            -- 
          begin -- 
            word_access_0_2439_start <= Xentry_2437_symbol; -- control passed to block
            Xentry_2440_symbol  <= word_access_0_2439_start; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/$entry
            cr_2442_symbol <= Xentry_2440_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/cr
            array_obj_ref_24_store_0_req_1 <= cr_2442_symbol; -- link to DP
            ca_2443_symbol <= array_obj_ref_24_store_0_ack_1; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/ca
            Xexit_2441_symbol <= ca_2443_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0/$exit
            word_access_0_2439_symbol <= Xexit_2441_symbol; -- control passed from block 
            -- 
          end Block; -- assign_stmt_26/array_obj_ref_24_complete/word_access/word_access_0
          Xexit_2438_symbol <= word_access_0_2439_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/word_access/$exit
          word_access_2436_symbol <= Xexit_2438_symbol; -- control passed from block 
          -- 
        end Block; -- assign_stmt_26/array_obj_ref_24_complete/word_access
        Xexit_2435_symbol <= word_access_2436_symbol; -- transition assign_stmt_26/array_obj_ref_24_complete/$exit
        array_obj_ref_24_complete_2433_symbol <= Xexit_2435_symbol; -- control passed from block 
        -- 
      end Block; -- assign_stmt_26/array_obj_ref_24_complete
      Xexit_2364_symbol <= assign_stmt_26_completed_x_x2366_symbol; -- transition assign_stmt_26/$exit
      assign_stmt_26_2362_symbol <= Xexit_2364_symbol; -- control passed from block 
      -- 
    end Block; -- assign_stmt_26
    Xexit_2361_symbol <= assign_stmt_26_2362_symbol; -- transition $exit
    fin  <=  '1' when Xexit_2361_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_24_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_24_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_word_address_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_24_word_offset_0 : std_logic_vector(0 downto 0);
    signal binary_21_wire : std_logic_vector(31 downto 0);
    signal binary_23_resized : std_logic_vector(0 downto 0);
    signal binary_23_scaled : std_logic_vector(0 downto 0);
    signal binary_23_wire : std_logic_vector(31 downto 0);
    signal expr_20_wire_constant : std_logic_vector(31 downto 0);
    signal expr_22_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_24_offset_scale_factor_0 <= "1";
    array_obj_ref_24_resized_base_address <= "0";
    array_obj_ref_24_word_offset_0 <= "0";
    expr_20_wire_constant <= "00000000000000000000000000000001";
    expr_22_wire_constant <= "00000000000000000000000000000000";
    array_obj_ref_24_index_0_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 1) -- 
      port map( din => binary_23_wire, dout => binary_23_resized, req => array_obj_ref_24_index_0_resize_req_0, ack => array_obj_ref_24_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_24_offset_inst: RegisterBase generic map(in_data_width => 1,out_data_width => 1) -- 
      port map( din => binary_23_scaled, dout => array_obj_ref_24_final_offset, req => array_obj_ref_24_offset_inst_req_0, ack => array_obj_ref_24_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_24_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_24_addr_0_ack_0 <= array_obj_ref_24_addr_0_req_0;
      aggregated_sig <= array_obj_ref_24_root_address;
      array_obj_ref_24_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_24_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_24_gather_scatter_ack_0 <= array_obj_ref_24_gather_scatter_req_0;
      aggregated_sig <= data;
      array_obj_ref_24_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_24_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_24_index_0_rename_ack_0 <= array_obj_ref_24_index_0_rename_req_0;
      aggregated_sig <= binary_23_resized;
      binary_23_scaled <= aggregated_sig(0 downto 0);
      --
    end Block;
    array_obj_ref_24_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      array_obj_ref_24_root_address_inst_ack_0 <= array_obj_ref_24_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_24_final_offset;
      array_obj_ref_24_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    -- shared split operator group (0) : binary_21_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= address;
      binary_21_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_21_inst_req_0,
          ackL => binary_21_inst_ack_0,
          reqR => binary_21_inst_req_1,
          ackR => binary_21_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_23_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_21_wire;
      binary_23_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000000",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_23_inst_req_0,
          ackL => binary_23_inst_ack_0,
          reqR => binary_23_inst_req_1,
          ackR => binary_23_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared store operator group (0) : array_obj_ref_24_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= array_obj_ref_24_store_0_req_0;
      array_obj_ref_24_store_0_ack_0 <= ackL(0);
      reqR(0) <= array_obj_ref_24_store_0_req_1;
      array_obj_ref_24_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_24_word_address_0;
      data_in <= array_obj_ref_24_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(0 downto 0),
          mdata => memory_space_0_sr_data(7 downto 0),
          mtag => memory_space_0_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity output_module is -- 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    foo_out_pipe_read_req : out  std_logic_vector(0 downto 0);
    foo_out_pipe_read_ack : in   std_logic_vector(0 downto 0);
    foo_out_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    output_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_data_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity output_module;
architecture Default of output_module is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_535_store_0_ack_1 : boolean;
  signal type_cast_528_inst_ack_0 : boolean;
  signal ptr_deref_535_gather_scatter_req_0 : boolean;
  signal type_cast_532_inst_req_0 : boolean;
  signal ptr_deref_540_load_0_req_1 : boolean;
  signal ptr_deref_535_gather_scatter_ack_0 : boolean;
  signal ptr_deref_571_gather_scatter_ack_0 : boolean;
  signal ptr_deref_540_gather_scatter_req_0 : boolean;
  signal ptr_deref_535_store_0_ack_0 : boolean;
  signal ptr_deref_571_load_0_ack_1 : boolean;
  signal ptr_deref_571_gather_scatter_req_0 : boolean;
  signal type_cast_532_inst_ack_0 : boolean;
  signal ptr_deref_540_load_0_req_0 : boolean;
  signal ptr_deref_540_load_0_ack_0 : boolean;
  signal ptr_deref_549_load_0_ack_1 : boolean;
  signal simple_obj_ref_556_inst_req_0 : boolean;
  signal simple_obj_ref_556_inst_ack_0 : boolean;
  signal ptr_deref_571_load_0_req_0 : boolean;
  signal type_cast_575_inst_ack_0 : boolean;
  signal type_cast_575_inst_req_0 : boolean;
  signal ptr_deref_549_gather_scatter_req_0 : boolean;
  signal ptr_deref_571_load_0_ack_0 : boolean;
  signal type_cast_558_inst_req_0 : boolean;
  signal type_cast_558_inst_ack_0 : boolean;
  signal ptr_deref_571_load_0_req_1 : boolean;
  signal ptr_deref_549_addr_0_req_0 : boolean;
  signal ptr_deref_549_addr_0_ack_0 : boolean;
  signal array_obj_ref_545_base_resize_ack_0 : boolean;
  signal ptr_deref_535_store_0_req_0 : boolean;
  signal ptr_deref_549_load_0_req_1 : boolean;
  signal array_obj_ref_545_base_resize_req_0 : boolean;
  signal ptr_deref_540_gather_scatter_ack_0 : boolean;
  signal ptr_deref_549_load_0_req_0 : boolean;
  signal ptr_deref_549_load_0_ack_0 : boolean;
  signal array_obj_ref_545_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_545_root_address_inst_req_1 : boolean;
  signal array_obj_ref_545_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_545_root_address_inst_req_0 : boolean;
  signal ptr_deref_549_gather_scatter_ack_0 : boolean;
  signal type_cast_528_inst_req_0 : boolean;
  signal simple_obj_ref_565_inst_ack_0 : boolean;
  signal ptr_deref_535_store_0_req_1 : boolean;
  signal array_obj_ref_545_final_reg_ack_0 : boolean;
  signal simple_obj_ref_565_inst_req_0 : boolean;
  signal ptr_deref_549_base_resize_req_0 : boolean;
  signal ptr_deref_549_base_resize_ack_0 : boolean;
  signal simple_obj_ref_527_inst_ack_0 : boolean;
  signal simple_obj_ref_527_inst_req_0 : boolean;
  signal ptr_deref_549_root_address_inst_req_0 : boolean;
  signal ptr_deref_549_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_545_final_reg_req_0 : boolean;
  signal ptr_deref_540_load_0_ack_1 : boolean;
  signal simple_obj_ref_582_inst_req_0 : boolean;
  signal simple_obj_ref_582_inst_ack_0 : boolean;
  signal type_cast_584_inst_req_0 : boolean;
  signal type_cast_584_inst_ack_0 : boolean;
  signal memory_space_17_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_17_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_17_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_17_lr_tag : std_logic_vector(1 downto 0);
  signal memory_space_17_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_17_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_17_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_17_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_17_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_17_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_17_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_17_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_17_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_17_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_17_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_17_sc_tag :  std_logic_vector(1 downto 0);
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  output_module_CP_2444: Block -- control-path 
    signal output_module_CP_2444_start: Boolean;
    signal Xentry_2445_symbol: Boolean;
    signal Xexit_2446_symbol: Boolean;
    signal branch_block_stmt_513_2447_symbol : Boolean;
    -- 
  begin -- 
    output_module_CP_2444_start <=  true when start = '1' else false; -- control passed to control-path.
    Xentry_2445_symbol  <= output_module_CP_2444_start; -- transition $entry
    branch_block_stmt_513_2447: Block -- branch_block_stmt_513 
      signal branch_block_stmt_513_2447_start: Boolean;
      signal Xentry_2448_symbol: Boolean;
      signal Xexit_2449_symbol: Boolean;
      signal branch_block_stmt_513_x_xentry_x_xx_x2450_symbol : Boolean;
      signal branch_block_stmt_513_x_xexit_x_xx_x2451_symbol : Boolean;
      signal assign_stmt_518_x_xentry_x_xx_x2452_symbol : Boolean;
      signal assign_stmt_518_x_xexit_x_xx_x2453_symbol : Boolean;
      signal bb_0_bb_1_2454_symbol : Boolean;
      signal merge_stmt_520_x_xexit_x_xx_x2455_symbol : Boolean;
      signal assign_stmt_525_x_xentry_x_xx_x2456_symbol : Boolean;
      signal assign_stmt_525_x_xexit_x_xx_x2457_symbol : Boolean;
      signal assign_stmt_529_x_xentry_x_xx_x2458_symbol : Boolean;
      signal assign_stmt_529_x_xexit_x_xx_x2459_symbol : Boolean;
      signal assign_stmt_533_to_assign_stmt_555_x_xentry_x_xx_x2460_symbol : Boolean;
      signal assign_stmt_533_to_assign_stmt_555_x_xexit_x_xx_x2461_symbol : Boolean;
      signal assign_stmt_559_x_xentry_x_xx_x2462_symbol : Boolean;
      signal assign_stmt_559_x_xexit_x_xx_x2463_symbol : Boolean;
      signal assign_stmt_564_x_xentry_x_xx_x2464_symbol : Boolean;
      signal assign_stmt_564_x_xexit_x_xx_x2465_symbol : Boolean;
      signal assign_stmt_568_x_xentry_x_xx_x2466_symbol : Boolean;
      signal assign_stmt_568_x_xexit_x_xx_x2467_symbol : Boolean;
      signal assign_stmt_572_to_assign_stmt_581_x_xentry_x_xx_x2468_symbol : Boolean;
      signal assign_stmt_572_to_assign_stmt_581_x_xexit_x_xx_x2469_symbol : Boolean;
      signal assign_stmt_585_x_xentry_x_xx_x2470_symbol : Boolean;
      signal assign_stmt_585_x_xexit_x_xx_x2471_symbol : Boolean;
      signal bb_1_bb_1_2472_symbol : Boolean;
      signal assign_stmt_518_2473_symbol : Boolean;
      signal assign_stmt_525_2476_symbol : Boolean;
      signal assign_stmt_529_2479_symbol : Boolean;
      signal assign_stmt_533_to_assign_stmt_555_2497_symbol : Boolean;
      signal assign_stmt_559_2646_symbol : Boolean;
      signal assign_stmt_564_2665_symbol : Boolean;
      signal assign_stmt_568_2668_symbol : Boolean;
      signal assign_stmt_572_to_assign_stmt_581_2679_symbol : Boolean;
      signal assign_stmt_585_2723_symbol : Boolean;
      signal bb_0_bb_1_PhiReq_2742_symbol : Boolean;
      signal bb_1_bb_1_PhiReq_2745_symbol : Boolean;
      signal merge_stmt_520_PhiReqMerge_2748_symbol : Boolean;
      signal merge_stmt_520_PhiAck_2749_symbol : Boolean;
      -- 
    begin -- 
      branch_block_stmt_513_2447_start <= Xentry_2445_symbol; -- control passed to block
      Xentry_2448_symbol  <= branch_block_stmt_513_2447_start; -- transition branch_block_stmt_513/$entry
      branch_block_stmt_513_x_xentry_x_xx_x2450_symbol  <=  Xentry_2448_symbol; -- place branch_block_stmt_513/branch_block_stmt_513__entry__ (optimized away) 
      branch_block_stmt_513_x_xexit_x_xx_x2451_symbol  <=   false ; -- place branch_block_stmt_513/branch_block_stmt_513__exit__ (optimized away) 
      assign_stmt_518_x_xentry_x_xx_x2452_symbol  <=  branch_block_stmt_513_x_xentry_x_xx_x2450_symbol; -- place branch_block_stmt_513/assign_stmt_518__entry__ (optimized away) 
      assign_stmt_518_x_xexit_x_xx_x2453_symbol  <=  assign_stmt_518_2473_symbol; -- place branch_block_stmt_513/assign_stmt_518__exit__ (optimized away) 
      bb_0_bb_1_2454_symbol  <=  assign_stmt_518_x_xexit_x_xx_x2453_symbol; -- place branch_block_stmt_513/bb_0_bb_1 (optimized away) 
      merge_stmt_520_x_xexit_x_xx_x2455_symbol  <=  merge_stmt_520_PhiAck_2749_symbol; -- place branch_block_stmt_513/merge_stmt_520__exit__ (optimized away) 
      assign_stmt_525_x_xentry_x_xx_x2456_symbol  <=  merge_stmt_520_x_xexit_x_xx_x2455_symbol; -- place branch_block_stmt_513/assign_stmt_525__entry__ (optimized away) 
      assign_stmt_525_x_xexit_x_xx_x2457_symbol  <=  assign_stmt_525_2476_symbol; -- place branch_block_stmt_513/assign_stmt_525__exit__ (optimized away) 
      assign_stmt_529_x_xentry_x_xx_x2458_symbol  <=  assign_stmt_525_x_xexit_x_xx_x2457_symbol; -- place branch_block_stmt_513/assign_stmt_529__entry__ (optimized away) 
      assign_stmt_529_x_xexit_x_xx_x2459_symbol  <=  assign_stmt_529_2479_symbol; -- place branch_block_stmt_513/assign_stmt_529__exit__ (optimized away) 
      assign_stmt_533_to_assign_stmt_555_x_xentry_x_xx_x2460_symbol  <=  assign_stmt_529_x_xexit_x_xx_x2459_symbol; -- place branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555__entry__ (optimized away) 
      assign_stmt_533_to_assign_stmt_555_x_xexit_x_xx_x2461_symbol  <=  assign_stmt_533_to_assign_stmt_555_2497_symbol; -- place branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555__exit__ (optimized away) 
      assign_stmt_559_x_xentry_x_xx_x2462_symbol  <=  assign_stmt_533_to_assign_stmt_555_x_xexit_x_xx_x2461_symbol; -- place branch_block_stmt_513/assign_stmt_559__entry__ (optimized away) 
      assign_stmt_559_x_xexit_x_xx_x2463_symbol  <=  assign_stmt_559_2646_symbol; -- place branch_block_stmt_513/assign_stmt_559__exit__ (optimized away) 
      assign_stmt_564_x_xentry_x_xx_x2464_symbol  <=  assign_stmt_559_x_xexit_x_xx_x2463_symbol; -- place branch_block_stmt_513/assign_stmt_564__entry__ (optimized away) 
      assign_stmt_564_x_xexit_x_xx_x2465_symbol  <=  assign_stmt_564_2665_symbol; -- place branch_block_stmt_513/assign_stmt_564__exit__ (optimized away) 
      assign_stmt_568_x_xentry_x_xx_x2466_symbol  <=  assign_stmt_564_x_xexit_x_xx_x2465_symbol; -- place branch_block_stmt_513/assign_stmt_568__entry__ (optimized away) 
      assign_stmt_568_x_xexit_x_xx_x2467_symbol  <=  assign_stmt_568_2668_symbol; -- place branch_block_stmt_513/assign_stmt_568__exit__ (optimized away) 
      assign_stmt_572_to_assign_stmt_581_x_xentry_x_xx_x2468_symbol  <=  assign_stmt_568_x_xexit_x_xx_x2467_symbol; -- place branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581__entry__ (optimized away) 
      assign_stmt_572_to_assign_stmt_581_x_xexit_x_xx_x2469_symbol  <=  assign_stmt_572_to_assign_stmt_581_2679_symbol; -- place branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581__exit__ (optimized away) 
      assign_stmt_585_x_xentry_x_xx_x2470_symbol  <=  assign_stmt_572_to_assign_stmt_581_x_xexit_x_xx_x2469_symbol; -- place branch_block_stmt_513/assign_stmt_585__entry__ (optimized away) 
      assign_stmt_585_x_xexit_x_xx_x2471_symbol  <=  assign_stmt_585_2723_symbol; -- place branch_block_stmt_513/assign_stmt_585__exit__ (optimized away) 
      bb_1_bb_1_2472_symbol  <=  assign_stmt_585_x_xexit_x_xx_x2471_symbol; -- place branch_block_stmt_513/bb_1_bb_1 (optimized away) 
      assign_stmt_518_2473: Block -- branch_block_stmt_513/assign_stmt_518 
        signal assign_stmt_518_2473_start: Boolean;
        signal Xentry_2474_symbol: Boolean;
        signal Xexit_2475_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_518_2473_start <= assign_stmt_518_x_xentry_x_xx_x2452_symbol; -- control passed to block
        Xentry_2474_symbol  <= assign_stmt_518_2473_start; -- transition branch_block_stmt_513/assign_stmt_518/$entry
        Xexit_2475_symbol <= Xentry_2474_symbol; -- transition branch_block_stmt_513/assign_stmt_518/$exit
        assign_stmt_518_2473_symbol <= Xexit_2475_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_518
      assign_stmt_525_2476: Block -- branch_block_stmt_513/assign_stmt_525 
        signal assign_stmt_525_2476_start: Boolean;
        signal Xentry_2477_symbol: Boolean;
        signal Xexit_2478_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_525_2476_start <= assign_stmt_525_x_xentry_x_xx_x2456_symbol; -- control passed to block
        Xentry_2477_symbol  <= assign_stmt_525_2476_start; -- transition branch_block_stmt_513/assign_stmt_525/$entry
        Xexit_2478_symbol <= Xentry_2477_symbol; -- transition branch_block_stmt_513/assign_stmt_525/$exit
        assign_stmt_525_2476_symbol <= Xexit_2478_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_525
      assign_stmt_529_2479: Block -- branch_block_stmt_513/assign_stmt_529 
        signal assign_stmt_529_2479_start: Boolean;
        signal Xentry_2480_symbol: Boolean;
        signal Xexit_2481_symbol: Boolean;
        signal assign_stmt_529_active_x_x2482_symbol : Boolean;
        signal assign_stmt_529_completed_x_x2483_symbol : Boolean;
        signal type_cast_528_active_x_x2484_symbol : Boolean;
        signal type_cast_528_trigger_x_x2485_symbol : Boolean;
        signal simple_obj_ref_527_trigger_x_x2486_symbol : Boolean;
        signal simple_obj_ref_527_complete_2487_symbol : Boolean;
        signal type_cast_528_complete_2492_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_529_2479_start <= assign_stmt_529_x_xentry_x_xx_x2458_symbol; -- control passed to block
        Xentry_2480_symbol  <= assign_stmt_529_2479_start; -- transition branch_block_stmt_513/assign_stmt_529/$entry
        assign_stmt_529_active_x_x2482_symbol <= type_cast_528_complete_2492_symbol; -- transition branch_block_stmt_513/assign_stmt_529/assign_stmt_529_active_
        assign_stmt_529_completed_x_x2483_symbol <= assign_stmt_529_active_x_x2482_symbol; -- transition branch_block_stmt_513/assign_stmt_529/assign_stmt_529_completed_
        type_cast_528_active_x_x2484_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_529/type_cast_528_active_ 
          signal type_cast_528_active_x_x2484_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_528_active_x_x2484_predecessors(0) <= type_cast_528_trigger_x_x2485_symbol;
          type_cast_528_active_x_x2484_predecessors(1) <= simple_obj_ref_527_complete_2487_symbol;
          type_cast_528_active_x_x2484_join: join -- 
            port map( -- 
              preds => type_cast_528_active_x_x2484_predecessors,
              symbol_out => type_cast_528_active_x_x2484_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_529/type_cast_528_active_
        type_cast_528_trigger_x_x2485_symbol <= Xentry_2480_symbol; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_trigger_
        simple_obj_ref_527_trigger_x_x2486_symbol <= Xentry_2480_symbol; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_trigger_
        simple_obj_ref_527_complete_2487: Block -- branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete 
          signal simple_obj_ref_527_complete_2487_start: Boolean;
          signal Xentry_2488_symbol: Boolean;
          signal Xexit_2489_symbol: Boolean;
          signal req_2490_symbol : Boolean;
          signal ack_2491_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_527_complete_2487_start <= simple_obj_ref_527_trigger_x_x2486_symbol; -- control passed to block
          Xentry_2488_symbol  <= simple_obj_ref_527_complete_2487_start; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/$entry
          req_2490_symbol <= Xentry_2488_symbol; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/req
          simple_obj_ref_527_inst_req_0 <= req_2490_symbol; -- link to DP
          ack_2491_symbol <= simple_obj_ref_527_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/ack
          Xexit_2489_symbol <= ack_2491_symbol; -- transition branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete/$exit
          simple_obj_ref_527_complete_2487_symbol <= Xexit_2489_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_529/simple_obj_ref_527_complete
        type_cast_528_complete_2492: Block -- branch_block_stmt_513/assign_stmt_529/type_cast_528_complete 
          signal type_cast_528_complete_2492_start: Boolean;
          signal Xentry_2493_symbol: Boolean;
          signal Xexit_2494_symbol: Boolean;
          signal req_2495_symbol : Boolean;
          signal ack_2496_symbol : Boolean;
          -- 
        begin -- 
          type_cast_528_complete_2492_start <= type_cast_528_active_x_x2484_symbol; -- control passed to block
          Xentry_2493_symbol  <= type_cast_528_complete_2492_start; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/$entry
          req_2495_symbol <= Xentry_2493_symbol; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/req
          type_cast_528_inst_req_0 <= req_2495_symbol; -- link to DP
          ack_2496_symbol <= type_cast_528_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/ack
          Xexit_2494_symbol <= ack_2496_symbol; -- transition branch_block_stmt_513/assign_stmt_529/type_cast_528_complete/$exit
          type_cast_528_complete_2492_symbol <= Xexit_2494_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_529/type_cast_528_complete
        Xexit_2481_symbol <= assign_stmt_529_completed_x_x2483_symbol; -- transition branch_block_stmt_513/assign_stmt_529/$exit
        assign_stmt_529_2479_symbol <= Xexit_2481_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_529
      assign_stmt_533_to_assign_stmt_555_2497: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555 
        signal assign_stmt_533_to_assign_stmt_555_2497_start: Boolean;
        signal Xentry_2498_symbol: Boolean;
        signal Xexit_2499_symbol: Boolean;
        signal assign_stmt_533_active_x_x2500_symbol : Boolean;
        signal assign_stmt_533_completed_x_x2501_symbol : Boolean;
        signal type_cast_532_active_x_x2502_symbol : Boolean;
        signal type_cast_532_trigger_x_x2503_symbol : Boolean;
        signal simple_obj_ref_531_complete_2504_symbol : Boolean;
        signal type_cast_532_complete_2505_symbol : Boolean;
        signal assign_stmt_537_active_x_x2510_symbol : Boolean;
        signal assign_stmt_537_completed_x_x2511_symbol : Boolean;
        signal simple_obj_ref_536_complete_2512_symbol : Boolean;
        signal ptr_deref_535_trigger_x_x2513_symbol : Boolean;
        signal ptr_deref_535_active_x_x2514_symbol : Boolean;
        signal ptr_deref_535_base_address_calculated_2515_symbol : Boolean;
        signal ptr_deref_535_root_address_calculated_2516_symbol : Boolean;
        signal ptr_deref_535_word_address_calculated_2517_symbol : Boolean;
        signal ptr_deref_535_request_2518_symbol : Boolean;
        signal ptr_deref_535_complete_2531_symbol : Boolean;
        signal assign_stmt_541_active_x_x2542_symbol : Boolean;
        signal assign_stmt_541_completed_x_x2543_symbol : Boolean;
        signal ptr_deref_540_trigger_x_x2544_symbol : Boolean;
        signal ptr_deref_540_active_x_x2545_symbol : Boolean;
        signal ptr_deref_540_base_address_calculated_2546_symbol : Boolean;
        signal ptr_deref_540_root_address_calculated_2547_symbol : Boolean;
        signal ptr_deref_540_word_address_calculated_2548_symbol : Boolean;
        signal ptr_deref_540_request_2549_symbol : Boolean;
        signal ptr_deref_540_complete_2560_symbol : Boolean;
        signal assign_stmt_546_active_x_x2573_symbol : Boolean;
        signal assign_stmt_546_completed_x_x2574_symbol : Boolean;
        signal array_obj_ref_545_trigger_x_x2575_symbol : Boolean;
        signal array_obj_ref_545_active_x_x2576_symbol : Boolean;
        signal array_obj_ref_545_base_address_calculated_2577_symbol : Boolean;
        signal array_obj_ref_545_root_address_calculated_2578_symbol : Boolean;
        signal array_obj_ref_545_base_address_resized_2579_symbol : Boolean;
        signal array_obj_ref_545_base_addr_resize_2580_symbol : Boolean;
        signal array_obj_ref_545_base_plus_offset_trigger_2585_symbol : Boolean;
        signal array_obj_ref_545_base_plus_offset_2586_symbol : Boolean;
        signal array_obj_ref_545_complete_2593_symbol : Boolean;
        signal assign_stmt_550_active_x_x2598_symbol : Boolean;
        signal assign_stmt_550_completed_x_x2599_symbol : Boolean;
        signal ptr_deref_549_trigger_x_x2600_symbol : Boolean;
        signal ptr_deref_549_active_x_x2601_symbol : Boolean;
        signal ptr_deref_549_base_address_calculated_2602_symbol : Boolean;
        signal simple_obj_ref_548_complete_2603_symbol : Boolean;
        signal ptr_deref_549_root_address_calculated_2604_symbol : Boolean;
        signal ptr_deref_549_word_address_calculated_2605_symbol : Boolean;
        signal ptr_deref_549_base_address_resized_2606_symbol : Boolean;
        signal ptr_deref_549_base_addr_resize_2607_symbol : Boolean;
        signal ptr_deref_549_base_plus_offset_2612_symbol : Boolean;
        signal ptr_deref_549_word_addrgen_2617_symbol : Boolean;
        signal ptr_deref_549_request_2622_symbol : Boolean;
        signal ptr_deref_549_complete_2633_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_533_to_assign_stmt_555_2497_start <= assign_stmt_533_to_assign_stmt_555_x_xentry_x_xx_x2460_symbol; -- control passed to block
        Xentry_2498_symbol  <= assign_stmt_533_to_assign_stmt_555_2497_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/$entry
        assign_stmt_533_active_x_x2500_symbol <= type_cast_532_complete_2505_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_533_active_
        assign_stmt_533_completed_x_x2501_symbol <= assign_stmt_533_active_x_x2500_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_533_completed_
        type_cast_532_active_x_x2502_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_active_ 
          signal type_cast_532_active_x_x2502_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_532_active_x_x2502_predecessors(0) <= type_cast_532_trigger_x_x2503_symbol;
          type_cast_532_active_x_x2502_predecessors(1) <= simple_obj_ref_531_complete_2504_symbol;
          type_cast_532_active_x_x2502_join: join -- 
            port map( -- 
              preds => type_cast_532_active_x_x2502_predecessors,
              symbol_out => type_cast_532_active_x_x2502_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_active_
        type_cast_532_trigger_x_x2503_symbol <= Xentry_2498_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_trigger_
        simple_obj_ref_531_complete_2504_symbol <= Xentry_2498_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/simple_obj_ref_531_complete
        type_cast_532_complete_2505: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete 
          signal type_cast_532_complete_2505_start: Boolean;
          signal Xentry_2506_symbol: Boolean;
          signal Xexit_2507_symbol: Boolean;
          signal req_2508_symbol : Boolean;
          signal ack_2509_symbol : Boolean;
          -- 
        begin -- 
          type_cast_532_complete_2505_start <= type_cast_532_active_x_x2502_symbol; -- control passed to block
          Xentry_2506_symbol  <= type_cast_532_complete_2505_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/$entry
          req_2508_symbol <= Xentry_2506_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/req
          type_cast_532_inst_req_0 <= req_2508_symbol; -- link to DP
          ack_2509_symbol <= type_cast_532_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/ack
          Xexit_2507_symbol <= ack_2509_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete/$exit
          type_cast_532_complete_2505_symbol <= Xexit_2507_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/type_cast_532_complete
        assign_stmt_537_active_x_x2510_symbol <= simple_obj_ref_536_complete_2512_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_537_active_
        assign_stmt_537_completed_x_x2511_symbol <= ptr_deref_535_complete_2531_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_537_completed_
        simple_obj_ref_536_complete_2512_symbol <= assign_stmt_533_completed_x_x2501_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/simple_obj_ref_536_complete
        ptr_deref_535_trigger_x_x2513_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_trigger_ 
          signal ptr_deref_535_trigger_x_x2513_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_535_trigger_x_x2513_predecessors(0) <= ptr_deref_535_word_address_calculated_2517_symbol;
          ptr_deref_535_trigger_x_x2513_predecessors(1) <= assign_stmt_537_active_x_x2510_symbol;
          ptr_deref_535_trigger_x_x2513_join: join -- 
            port map( -- 
              preds => ptr_deref_535_trigger_x_x2513_predecessors,
              symbol_out => ptr_deref_535_trigger_x_x2513_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_trigger_
        ptr_deref_535_active_x_x2514_symbol <= ptr_deref_535_request_2518_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_active_
        ptr_deref_535_base_address_calculated_2515_symbol <= Xentry_2498_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_base_address_calculated
        ptr_deref_535_root_address_calculated_2516_symbol <= Xentry_2498_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_root_address_calculated
        ptr_deref_535_word_address_calculated_2517_symbol <= ptr_deref_535_root_address_calculated_2516_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_word_address_calculated
        ptr_deref_535_request_2518: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request 
          signal ptr_deref_535_request_2518_start: Boolean;
          signal Xentry_2519_symbol: Boolean;
          signal Xexit_2520_symbol: Boolean;
          signal split_req_2521_symbol : Boolean;
          signal split_ack_2522_symbol : Boolean;
          signal word_access_2523_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_535_request_2518_start <= ptr_deref_535_trigger_x_x2513_symbol; -- control passed to block
          Xentry_2519_symbol  <= ptr_deref_535_request_2518_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/$entry
          split_req_2521_symbol <= Xentry_2519_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/split_req
          ptr_deref_535_gather_scatter_req_0 <= split_req_2521_symbol; -- link to DP
          split_ack_2522_symbol <= ptr_deref_535_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/split_ack
          word_access_2523: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access 
            signal word_access_2523_start: Boolean;
            signal Xentry_2524_symbol: Boolean;
            signal Xexit_2525_symbol: Boolean;
            signal word_access_0_2526_symbol : Boolean;
            -- 
          begin -- 
            word_access_2523_start <= split_ack_2522_symbol; -- control passed to block
            Xentry_2524_symbol  <= word_access_2523_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/$entry
            word_access_0_2526: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0 
              signal word_access_0_2526_start: Boolean;
              signal Xentry_2527_symbol: Boolean;
              signal Xexit_2528_symbol: Boolean;
              signal rr_2529_symbol : Boolean;
              signal ra_2530_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2526_start <= Xentry_2524_symbol; -- control passed to block
              Xentry_2527_symbol  <= word_access_0_2526_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/$entry
              rr_2529_symbol <= Xentry_2527_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/rr
              ptr_deref_535_store_0_req_0 <= rr_2529_symbol; -- link to DP
              ra_2530_symbol <= ptr_deref_535_store_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/ra
              Xexit_2528_symbol <= ra_2530_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0/$exit
              word_access_0_2526_symbol <= Xexit_2528_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/word_access_0
            Xexit_2525_symbol <= word_access_0_2526_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access/$exit
            word_access_2523_symbol <= Xexit_2525_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/word_access
          Xexit_2520_symbol <= word_access_2523_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request/$exit
          ptr_deref_535_request_2518_symbol <= Xexit_2520_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_request
        ptr_deref_535_complete_2531: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete 
          signal ptr_deref_535_complete_2531_start: Boolean;
          signal Xentry_2532_symbol: Boolean;
          signal Xexit_2533_symbol: Boolean;
          signal word_access_2534_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_535_complete_2531_start <= ptr_deref_535_active_x_x2514_symbol; -- control passed to block
          Xentry_2532_symbol  <= ptr_deref_535_complete_2531_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/$entry
          word_access_2534: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access 
            signal word_access_2534_start: Boolean;
            signal Xentry_2535_symbol: Boolean;
            signal Xexit_2536_symbol: Boolean;
            signal word_access_0_2537_symbol : Boolean;
            -- 
          begin -- 
            word_access_2534_start <= Xentry_2532_symbol; -- control passed to block
            Xentry_2535_symbol  <= word_access_2534_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/$entry
            word_access_0_2537: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0 
              signal word_access_0_2537_start: Boolean;
              signal Xentry_2538_symbol: Boolean;
              signal Xexit_2539_symbol: Boolean;
              signal cr_2540_symbol : Boolean;
              signal ca_2541_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2537_start <= Xentry_2535_symbol; -- control passed to block
              Xentry_2538_symbol  <= word_access_0_2537_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/$entry
              cr_2540_symbol <= Xentry_2538_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/cr
              ptr_deref_535_store_0_req_1 <= cr_2540_symbol; -- link to DP
              ca_2541_symbol <= ptr_deref_535_store_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/ca
              Xexit_2539_symbol <= ca_2541_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0/$exit
              word_access_0_2537_symbol <= Xexit_2539_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/word_access_0
            Xexit_2536_symbol <= word_access_0_2537_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access/$exit
            word_access_2534_symbol <= Xexit_2536_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/word_access
          Xexit_2533_symbol <= word_access_2534_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete/$exit
          ptr_deref_535_complete_2531_symbol <= Xexit_2533_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_535_complete
        assign_stmt_541_active_x_x2542_symbol <= ptr_deref_540_complete_2560_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_541_active_
        assign_stmt_541_completed_x_x2543_symbol <= assign_stmt_541_active_x_x2542_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_541_completed_
        ptr_deref_540_trigger_x_x2544_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_trigger_ 
          signal ptr_deref_540_trigger_x_x2544_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_540_trigger_x_x2544_predecessors(0) <= ptr_deref_540_word_address_calculated_2548_symbol;
          ptr_deref_540_trigger_x_x2544_predecessors(1) <= ptr_deref_535_active_x_x2514_symbol;
          ptr_deref_540_trigger_x_x2544_join: join -- 
            port map( -- 
              preds => ptr_deref_540_trigger_x_x2544_predecessors,
              symbol_out => ptr_deref_540_trigger_x_x2544_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_trigger_
        ptr_deref_540_active_x_x2545_symbol <= ptr_deref_540_request_2549_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_active_
        ptr_deref_540_base_address_calculated_2546_symbol <= Xentry_2498_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_base_address_calculated
        ptr_deref_540_root_address_calculated_2547_symbol <= Xentry_2498_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_root_address_calculated
        ptr_deref_540_word_address_calculated_2548_symbol <= ptr_deref_540_root_address_calculated_2547_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_word_address_calculated
        ptr_deref_540_request_2549: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request 
          signal ptr_deref_540_request_2549_start: Boolean;
          signal Xentry_2550_symbol: Boolean;
          signal Xexit_2551_symbol: Boolean;
          signal word_access_2552_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_540_request_2549_start <= ptr_deref_540_trigger_x_x2544_symbol; -- control passed to block
          Xentry_2550_symbol  <= ptr_deref_540_request_2549_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/$entry
          word_access_2552: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access 
            signal word_access_2552_start: Boolean;
            signal Xentry_2553_symbol: Boolean;
            signal Xexit_2554_symbol: Boolean;
            signal word_access_0_2555_symbol : Boolean;
            -- 
          begin -- 
            word_access_2552_start <= Xentry_2550_symbol; -- control passed to block
            Xentry_2553_symbol  <= word_access_2552_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/$entry
            word_access_0_2555: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0 
              signal word_access_0_2555_start: Boolean;
              signal Xentry_2556_symbol: Boolean;
              signal Xexit_2557_symbol: Boolean;
              signal rr_2558_symbol : Boolean;
              signal ra_2559_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2555_start <= Xentry_2553_symbol; -- control passed to block
              Xentry_2556_symbol  <= word_access_0_2555_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/$entry
              rr_2558_symbol <= Xentry_2556_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/rr
              ptr_deref_540_load_0_req_0 <= rr_2558_symbol; -- link to DP
              ra_2559_symbol <= ptr_deref_540_load_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/ra
              Xexit_2557_symbol <= ra_2559_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0/$exit
              word_access_0_2555_symbol <= Xexit_2557_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/word_access_0
            Xexit_2554_symbol <= word_access_0_2555_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access/$exit
            word_access_2552_symbol <= Xexit_2554_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/word_access
          Xexit_2551_symbol <= word_access_2552_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request/$exit
          ptr_deref_540_request_2549_symbol <= Xexit_2551_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_request
        ptr_deref_540_complete_2560: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete 
          signal ptr_deref_540_complete_2560_start: Boolean;
          signal Xentry_2561_symbol: Boolean;
          signal Xexit_2562_symbol: Boolean;
          signal word_access_2563_symbol : Boolean;
          signal merge_req_2571_symbol : Boolean;
          signal merge_ack_2572_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_540_complete_2560_start <= ptr_deref_540_active_x_x2545_symbol; -- control passed to block
          Xentry_2561_symbol  <= ptr_deref_540_complete_2560_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/$entry
          word_access_2563: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access 
            signal word_access_2563_start: Boolean;
            signal Xentry_2564_symbol: Boolean;
            signal Xexit_2565_symbol: Boolean;
            signal word_access_0_2566_symbol : Boolean;
            -- 
          begin -- 
            word_access_2563_start <= Xentry_2561_symbol; -- control passed to block
            Xentry_2564_symbol  <= word_access_2563_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/$entry
            word_access_0_2566: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0 
              signal word_access_0_2566_start: Boolean;
              signal Xentry_2567_symbol: Boolean;
              signal Xexit_2568_symbol: Boolean;
              signal cr_2569_symbol : Boolean;
              signal ca_2570_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2566_start <= Xentry_2564_symbol; -- control passed to block
              Xentry_2567_symbol  <= word_access_0_2566_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/$entry
              cr_2569_symbol <= Xentry_2567_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/cr
              ptr_deref_540_load_0_req_1 <= cr_2569_symbol; -- link to DP
              ca_2570_symbol <= ptr_deref_540_load_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/ca
              Xexit_2568_symbol <= ca_2570_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0/$exit
              word_access_0_2566_symbol <= Xexit_2568_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/word_access_0
            Xexit_2565_symbol <= word_access_0_2566_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access/$exit
            word_access_2563_symbol <= Xexit_2565_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/word_access
          merge_req_2571_symbol <= word_access_2563_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/merge_req
          ptr_deref_540_gather_scatter_req_0 <= merge_req_2571_symbol; -- link to DP
          merge_ack_2572_symbol <= ptr_deref_540_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/merge_ack
          Xexit_2562_symbol <= merge_ack_2572_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete/$exit
          ptr_deref_540_complete_2560_symbol <= Xexit_2562_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_540_complete
        assign_stmt_546_active_x_x2573_symbol <= array_obj_ref_545_complete_2593_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_546_active_
        assign_stmt_546_completed_x_x2574_symbol <= assign_stmt_546_active_x_x2573_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_546_completed_
        array_obj_ref_545_trigger_x_x2575_symbol <= Xentry_2498_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_trigger_
        array_obj_ref_545_active_x_x2576_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_active_ 
          signal array_obj_ref_545_active_x_x2576_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          array_obj_ref_545_active_x_x2576_predecessors(0) <= array_obj_ref_545_trigger_x_x2575_symbol;
          array_obj_ref_545_active_x_x2576_predecessors(1) <= array_obj_ref_545_root_address_calculated_2578_symbol;
          array_obj_ref_545_active_x_x2576_join: join -- 
            port map( -- 
              preds => array_obj_ref_545_active_x_x2576_predecessors,
              symbol_out => array_obj_ref_545_active_x_x2576_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_active_
        array_obj_ref_545_base_address_calculated_2577_symbol <= assign_stmt_541_completed_x_x2543_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_address_calculated
        array_obj_ref_545_root_address_calculated_2578_symbol <= array_obj_ref_545_base_plus_offset_2586_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_root_address_calculated
        array_obj_ref_545_base_address_resized_2579_symbol <= array_obj_ref_545_base_addr_resize_2580_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_address_resized
        array_obj_ref_545_base_addr_resize_2580: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize 
          signal array_obj_ref_545_base_addr_resize_2580_start: Boolean;
          signal Xentry_2581_symbol: Boolean;
          signal Xexit_2582_symbol: Boolean;
          signal base_resize_req_2583_symbol : Boolean;
          signal base_resize_ack_2584_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_545_base_addr_resize_2580_start <= array_obj_ref_545_base_address_calculated_2577_symbol; -- control passed to block
          Xentry_2581_symbol  <= array_obj_ref_545_base_addr_resize_2580_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/$entry
          base_resize_req_2583_symbol <= Xentry_2581_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/base_resize_req
          array_obj_ref_545_base_resize_req_0 <= base_resize_req_2583_symbol; -- link to DP
          base_resize_ack_2584_symbol <= array_obj_ref_545_base_resize_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/base_resize_ack
          Xexit_2582_symbol <= base_resize_ack_2584_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize/$exit
          array_obj_ref_545_base_addr_resize_2580_symbol <= Xexit_2582_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_addr_resize
        array_obj_ref_545_base_plus_offset_trigger_2585_symbol <= array_obj_ref_545_base_address_resized_2579_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset_trigger
        array_obj_ref_545_base_plus_offset_2586: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset 
          signal array_obj_ref_545_base_plus_offset_2586_start: Boolean;
          signal Xentry_2587_symbol: Boolean;
          signal Xexit_2588_symbol: Boolean;
          signal plus_base_rr_2589_symbol : Boolean;
          signal plus_base_ra_2590_symbol : Boolean;
          signal plus_base_cr_2591_symbol : Boolean;
          signal plus_base_ca_2592_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_545_base_plus_offset_2586_start <= array_obj_ref_545_base_plus_offset_trigger_2585_symbol; -- control passed to block
          Xentry_2587_symbol  <= array_obj_ref_545_base_plus_offset_2586_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/$entry
          plus_base_rr_2589_symbol <= Xentry_2587_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_rr
          array_obj_ref_545_root_address_inst_req_0 <= plus_base_rr_2589_symbol; -- link to DP
          plus_base_ra_2590_symbol <= array_obj_ref_545_root_address_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_ra
          plus_base_cr_2591_symbol <= plus_base_ra_2590_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_cr
          array_obj_ref_545_root_address_inst_req_1 <= plus_base_cr_2591_symbol; -- link to DP
          plus_base_ca_2592_symbol <= array_obj_ref_545_root_address_inst_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/plus_base_ca
          Xexit_2588_symbol <= plus_base_ca_2592_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset/$exit
          array_obj_ref_545_base_plus_offset_2586_symbol <= Xexit_2588_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_base_plus_offset
        array_obj_ref_545_complete_2593: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete 
          signal array_obj_ref_545_complete_2593_start: Boolean;
          signal Xentry_2594_symbol: Boolean;
          signal Xexit_2595_symbol: Boolean;
          signal final_reg_req_2596_symbol : Boolean;
          signal final_reg_ack_2597_symbol : Boolean;
          -- 
        begin -- 
          array_obj_ref_545_complete_2593_start <= array_obj_ref_545_active_x_x2576_symbol; -- control passed to block
          Xentry_2594_symbol  <= array_obj_ref_545_complete_2593_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/$entry
          final_reg_req_2596_symbol <= Xentry_2594_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/final_reg_req
          array_obj_ref_545_final_reg_req_0 <= final_reg_req_2596_symbol; -- link to DP
          final_reg_ack_2597_symbol <= array_obj_ref_545_final_reg_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/final_reg_ack
          Xexit_2595_symbol <= final_reg_ack_2597_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete/$exit
          array_obj_ref_545_complete_2593_symbol <= Xexit_2595_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/array_obj_ref_545_complete
        assign_stmt_550_active_x_x2598_symbol <= ptr_deref_549_complete_2633_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_550_active_
        assign_stmt_550_completed_x_x2599_symbol <= assign_stmt_550_active_x_x2598_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/assign_stmt_550_completed_
        ptr_deref_549_trigger_x_x2600_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_trigger_ 
          signal ptr_deref_549_trigger_x_x2600_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          ptr_deref_549_trigger_x_x2600_predecessors(0) <= ptr_deref_549_word_address_calculated_2605_symbol;
          ptr_deref_549_trigger_x_x2600_predecessors(1) <= ptr_deref_549_base_address_calculated_2602_symbol;
          ptr_deref_549_trigger_x_x2600_join: join -- 
            port map( -- 
              preds => ptr_deref_549_trigger_x_x2600_predecessors,
              symbol_out => ptr_deref_549_trigger_x_x2600_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_trigger_
        ptr_deref_549_active_x_x2601_symbol <= ptr_deref_549_request_2622_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_active_
        ptr_deref_549_base_address_calculated_2602_symbol <= simple_obj_ref_548_complete_2603_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_address_calculated
        simple_obj_ref_548_complete_2603_symbol <= assign_stmt_546_completed_x_x2574_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/simple_obj_ref_548_complete
        ptr_deref_549_root_address_calculated_2604_symbol <= ptr_deref_549_base_plus_offset_2612_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_root_address_calculated
        ptr_deref_549_word_address_calculated_2605_symbol <= ptr_deref_549_word_addrgen_2617_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_address_calculated
        ptr_deref_549_base_address_resized_2606_symbol <= ptr_deref_549_base_addr_resize_2607_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_address_resized
        ptr_deref_549_base_addr_resize_2607: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize 
          signal ptr_deref_549_base_addr_resize_2607_start: Boolean;
          signal Xentry_2608_symbol: Boolean;
          signal Xexit_2609_symbol: Boolean;
          signal base_resize_req_2610_symbol : Boolean;
          signal base_resize_ack_2611_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_base_addr_resize_2607_start <= ptr_deref_549_base_address_calculated_2602_symbol; -- control passed to block
          Xentry_2608_symbol  <= ptr_deref_549_base_addr_resize_2607_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/$entry
          base_resize_req_2610_symbol <= Xentry_2608_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/base_resize_req
          ptr_deref_549_base_resize_req_0 <= base_resize_req_2610_symbol; -- link to DP
          base_resize_ack_2611_symbol <= ptr_deref_549_base_resize_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/base_resize_ack
          Xexit_2609_symbol <= base_resize_ack_2611_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize/$exit
          ptr_deref_549_base_addr_resize_2607_symbol <= Xexit_2609_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_addr_resize
        ptr_deref_549_base_plus_offset_2612: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset 
          signal ptr_deref_549_base_plus_offset_2612_start: Boolean;
          signal Xentry_2613_symbol: Boolean;
          signal Xexit_2614_symbol: Boolean;
          signal sum_rename_req_2615_symbol : Boolean;
          signal sum_rename_ack_2616_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_base_plus_offset_2612_start <= ptr_deref_549_base_address_resized_2606_symbol; -- control passed to block
          Xentry_2613_symbol  <= ptr_deref_549_base_plus_offset_2612_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/$entry
          sum_rename_req_2615_symbol <= Xentry_2613_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/sum_rename_req
          ptr_deref_549_root_address_inst_req_0 <= sum_rename_req_2615_symbol; -- link to DP
          sum_rename_ack_2616_symbol <= ptr_deref_549_root_address_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/sum_rename_ack
          Xexit_2614_symbol <= sum_rename_ack_2616_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset/$exit
          ptr_deref_549_base_plus_offset_2612_symbol <= Xexit_2614_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_base_plus_offset
        ptr_deref_549_word_addrgen_2617: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen 
          signal ptr_deref_549_word_addrgen_2617_start: Boolean;
          signal Xentry_2618_symbol: Boolean;
          signal Xexit_2619_symbol: Boolean;
          signal root_rename_req_2620_symbol : Boolean;
          signal root_rename_ack_2621_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_word_addrgen_2617_start <= ptr_deref_549_root_address_calculated_2604_symbol; -- control passed to block
          Xentry_2618_symbol  <= ptr_deref_549_word_addrgen_2617_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/$entry
          root_rename_req_2620_symbol <= Xentry_2618_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/root_rename_req
          ptr_deref_549_addr_0_req_0 <= root_rename_req_2620_symbol; -- link to DP
          root_rename_ack_2621_symbol <= ptr_deref_549_addr_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/root_rename_ack
          Xexit_2619_symbol <= root_rename_ack_2621_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen/$exit
          ptr_deref_549_word_addrgen_2617_symbol <= Xexit_2619_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_word_addrgen
        ptr_deref_549_request_2622: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request 
          signal ptr_deref_549_request_2622_start: Boolean;
          signal Xentry_2623_symbol: Boolean;
          signal Xexit_2624_symbol: Boolean;
          signal word_access_2625_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_request_2622_start <= ptr_deref_549_trigger_x_x2600_symbol; -- control passed to block
          Xentry_2623_symbol  <= ptr_deref_549_request_2622_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/$entry
          word_access_2625: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access 
            signal word_access_2625_start: Boolean;
            signal Xentry_2626_symbol: Boolean;
            signal Xexit_2627_symbol: Boolean;
            signal word_access_0_2628_symbol : Boolean;
            -- 
          begin -- 
            word_access_2625_start <= Xentry_2623_symbol; -- control passed to block
            Xentry_2626_symbol  <= word_access_2625_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/$entry
            word_access_0_2628: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0 
              signal word_access_0_2628_start: Boolean;
              signal Xentry_2629_symbol: Boolean;
              signal Xexit_2630_symbol: Boolean;
              signal rr_2631_symbol : Boolean;
              signal ra_2632_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2628_start <= Xentry_2626_symbol; -- control passed to block
              Xentry_2629_symbol  <= word_access_0_2628_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/$entry
              rr_2631_symbol <= Xentry_2629_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/rr
              ptr_deref_549_load_0_req_0 <= rr_2631_symbol; -- link to DP
              ra_2632_symbol <= ptr_deref_549_load_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/ra
              Xexit_2630_symbol <= ra_2632_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0/$exit
              word_access_0_2628_symbol <= Xexit_2630_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/word_access_0
            Xexit_2627_symbol <= word_access_0_2628_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access/$exit
            word_access_2625_symbol <= Xexit_2627_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/word_access
          Xexit_2624_symbol <= word_access_2625_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request/$exit
          ptr_deref_549_request_2622_symbol <= Xexit_2624_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_request
        ptr_deref_549_complete_2633: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete 
          signal ptr_deref_549_complete_2633_start: Boolean;
          signal Xentry_2634_symbol: Boolean;
          signal Xexit_2635_symbol: Boolean;
          signal word_access_2636_symbol : Boolean;
          signal merge_req_2644_symbol : Boolean;
          signal merge_ack_2645_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_549_complete_2633_start <= ptr_deref_549_active_x_x2601_symbol; -- control passed to block
          Xentry_2634_symbol  <= ptr_deref_549_complete_2633_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/$entry
          word_access_2636: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access 
            signal word_access_2636_start: Boolean;
            signal Xentry_2637_symbol: Boolean;
            signal Xexit_2638_symbol: Boolean;
            signal word_access_0_2639_symbol : Boolean;
            -- 
          begin -- 
            word_access_2636_start <= Xentry_2634_symbol; -- control passed to block
            Xentry_2637_symbol  <= word_access_2636_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/$entry
            word_access_0_2639: Block -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0 
              signal word_access_0_2639_start: Boolean;
              signal Xentry_2640_symbol: Boolean;
              signal Xexit_2641_symbol: Boolean;
              signal cr_2642_symbol : Boolean;
              signal ca_2643_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2639_start <= Xentry_2637_symbol; -- control passed to block
              Xentry_2640_symbol  <= word_access_0_2639_start; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/$entry
              cr_2642_symbol <= Xentry_2640_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/cr
              ptr_deref_549_load_0_req_1 <= cr_2642_symbol; -- link to DP
              ca_2643_symbol <= ptr_deref_549_load_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/ca
              Xexit_2641_symbol <= ca_2643_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0/$exit
              word_access_0_2639_symbol <= Xexit_2641_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/word_access_0
            Xexit_2638_symbol <= word_access_0_2639_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access/$exit
            word_access_2636_symbol <= Xexit_2638_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/word_access
          merge_req_2644_symbol <= word_access_2636_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/merge_req
          ptr_deref_549_gather_scatter_req_0 <= merge_req_2644_symbol; -- link to DP
          merge_ack_2645_symbol <= ptr_deref_549_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/merge_ack
          Xexit_2635_symbol <= merge_ack_2645_symbol; -- transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete/$exit
          ptr_deref_549_complete_2633_symbol <= Xexit_2635_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/ptr_deref_549_complete
        Xexit_2499_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/$exit 
          signal Xexit_2499_predecessors: BooleanArray(3 downto 0);
          -- 
        begin -- 
          Xexit_2499_predecessors(0) <= assign_stmt_537_completed_x_x2511_symbol;
          Xexit_2499_predecessors(1) <= ptr_deref_535_base_address_calculated_2515_symbol;
          Xexit_2499_predecessors(2) <= ptr_deref_540_base_address_calculated_2546_symbol;
          Xexit_2499_predecessors(3) <= assign_stmt_550_completed_x_x2599_symbol;
          Xexit_2499_join: join -- 
            port map( -- 
              preds => Xexit_2499_predecessors,
              symbol_out => Xexit_2499_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555/$exit
        assign_stmt_533_to_assign_stmt_555_2497_symbol <= Xexit_2499_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_533_to_assign_stmt_555
      assign_stmt_559_2646: Block -- branch_block_stmt_513/assign_stmt_559 
        signal assign_stmt_559_2646_start: Boolean;
        signal Xentry_2647_symbol: Boolean;
        signal Xexit_2648_symbol: Boolean;
        signal assign_stmt_559_active_x_x2649_symbol : Boolean;
        signal assign_stmt_559_completed_x_x2650_symbol : Boolean;
        signal type_cast_558_active_x_x2651_symbol : Boolean;
        signal type_cast_558_trigger_x_x2652_symbol : Boolean;
        signal simple_obj_ref_557_complete_2653_symbol : Boolean;
        signal type_cast_558_complete_2654_symbol : Boolean;
        signal simple_obj_ref_556_trigger_x_x2659_symbol : Boolean;
        signal simple_obj_ref_556_complete_2660_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_559_2646_start <= assign_stmt_559_x_xentry_x_xx_x2462_symbol; -- control passed to block
        Xentry_2647_symbol  <= assign_stmt_559_2646_start; -- transition branch_block_stmt_513/assign_stmt_559/$entry
        assign_stmt_559_active_x_x2649_symbol <= type_cast_558_complete_2654_symbol; -- transition branch_block_stmt_513/assign_stmt_559/assign_stmt_559_active_
        assign_stmt_559_completed_x_x2650_symbol <= simple_obj_ref_556_complete_2660_symbol; -- transition branch_block_stmt_513/assign_stmt_559/assign_stmt_559_completed_
        type_cast_558_active_x_x2651_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_559/type_cast_558_active_ 
          signal type_cast_558_active_x_x2651_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_558_active_x_x2651_predecessors(0) <= type_cast_558_trigger_x_x2652_symbol;
          type_cast_558_active_x_x2651_predecessors(1) <= simple_obj_ref_557_complete_2653_symbol;
          type_cast_558_active_x_x2651_join: join -- 
            port map( -- 
              preds => type_cast_558_active_x_x2651_predecessors,
              symbol_out => type_cast_558_active_x_x2651_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_559/type_cast_558_active_
        type_cast_558_trigger_x_x2652_symbol <= Xentry_2647_symbol; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_trigger_
        simple_obj_ref_557_complete_2653_symbol <= Xentry_2647_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_557_complete
        type_cast_558_complete_2654: Block -- branch_block_stmt_513/assign_stmt_559/type_cast_558_complete 
          signal type_cast_558_complete_2654_start: Boolean;
          signal Xentry_2655_symbol: Boolean;
          signal Xexit_2656_symbol: Boolean;
          signal req_2657_symbol : Boolean;
          signal ack_2658_symbol : Boolean;
          -- 
        begin -- 
          type_cast_558_complete_2654_start <= type_cast_558_active_x_x2651_symbol; -- control passed to block
          Xentry_2655_symbol  <= type_cast_558_complete_2654_start; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/$entry
          req_2657_symbol <= Xentry_2655_symbol; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/req
          type_cast_558_inst_req_0 <= req_2657_symbol; -- link to DP
          ack_2658_symbol <= type_cast_558_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/ack
          Xexit_2656_symbol <= ack_2658_symbol; -- transition branch_block_stmt_513/assign_stmt_559/type_cast_558_complete/$exit
          type_cast_558_complete_2654_symbol <= Xexit_2656_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_559/type_cast_558_complete
        simple_obj_ref_556_trigger_x_x2659_symbol <= assign_stmt_559_active_x_x2649_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_trigger_
        simple_obj_ref_556_complete_2660: Block -- branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete 
          signal simple_obj_ref_556_complete_2660_start: Boolean;
          signal Xentry_2661_symbol: Boolean;
          signal Xexit_2662_symbol: Boolean;
          signal pipe_wreq_2663_symbol : Boolean;
          signal pipe_wack_2664_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_556_complete_2660_start <= simple_obj_ref_556_trigger_x_x2659_symbol; -- control passed to block
          Xentry_2661_symbol  <= simple_obj_ref_556_complete_2660_start; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/$entry
          pipe_wreq_2663_symbol <= Xentry_2661_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/pipe_wreq
          simple_obj_ref_556_inst_req_0 <= pipe_wreq_2663_symbol; -- link to DP
          pipe_wack_2664_symbol <= simple_obj_ref_556_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/pipe_wack
          Xexit_2662_symbol <= pipe_wack_2664_symbol; -- transition branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete/$exit
          simple_obj_ref_556_complete_2660_symbol <= Xexit_2662_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_559/simple_obj_ref_556_complete
        Xexit_2648_symbol <= assign_stmt_559_completed_x_x2650_symbol; -- transition branch_block_stmt_513/assign_stmt_559/$exit
        assign_stmt_559_2646_symbol <= Xexit_2648_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_559
      assign_stmt_564_2665: Block -- branch_block_stmt_513/assign_stmt_564 
        signal assign_stmt_564_2665_start: Boolean;
        signal Xentry_2666_symbol: Boolean;
        signal Xexit_2667_symbol: Boolean;
        -- 
      begin -- 
        assign_stmt_564_2665_start <= assign_stmt_564_x_xentry_x_xx_x2464_symbol; -- control passed to block
        Xentry_2666_symbol  <= assign_stmt_564_2665_start; -- transition branch_block_stmt_513/assign_stmt_564/$entry
        Xexit_2667_symbol <= Xentry_2666_symbol; -- transition branch_block_stmt_513/assign_stmt_564/$exit
        assign_stmt_564_2665_symbol <= Xexit_2667_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_564
      assign_stmt_568_2668: Block -- branch_block_stmt_513/assign_stmt_568 
        signal assign_stmt_568_2668_start: Boolean;
        signal Xentry_2669_symbol: Boolean;
        signal Xexit_2670_symbol: Boolean;
        signal assign_stmt_568_active_x_x2671_symbol : Boolean;
        signal assign_stmt_568_completed_x_x2672_symbol : Boolean;
        signal simple_obj_ref_565_trigger_x_x2673_symbol : Boolean;
        signal simple_obj_ref_565_complete_2674_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_568_2668_start <= assign_stmt_568_x_xentry_x_xx_x2466_symbol; -- control passed to block
        Xentry_2669_symbol  <= assign_stmt_568_2668_start; -- transition branch_block_stmt_513/assign_stmt_568/$entry
        assign_stmt_568_active_x_x2671_symbol <= Xentry_2669_symbol; -- transition branch_block_stmt_513/assign_stmt_568/assign_stmt_568_active_
        assign_stmt_568_completed_x_x2672_symbol <= simple_obj_ref_565_complete_2674_symbol; -- transition branch_block_stmt_513/assign_stmt_568/assign_stmt_568_completed_
        simple_obj_ref_565_trigger_x_x2673_symbol <= assign_stmt_568_active_x_x2671_symbol; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_trigger_
        simple_obj_ref_565_complete_2674: Block -- branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete 
          signal simple_obj_ref_565_complete_2674_start: Boolean;
          signal Xentry_2675_symbol: Boolean;
          signal Xexit_2676_symbol: Boolean;
          signal pipe_wreq_2677_symbol : Boolean;
          signal pipe_wack_2678_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_565_complete_2674_start <= simple_obj_ref_565_trigger_x_x2673_symbol; -- control passed to block
          Xentry_2675_symbol  <= simple_obj_ref_565_complete_2674_start; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/$entry
          pipe_wreq_2677_symbol <= Xentry_2675_symbol; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/pipe_wreq
          simple_obj_ref_565_inst_req_0 <= pipe_wreq_2677_symbol; -- link to DP
          pipe_wack_2678_symbol <= simple_obj_ref_565_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/pipe_wack
          Xexit_2676_symbol <= pipe_wack_2678_symbol; -- transition branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete/$exit
          simple_obj_ref_565_complete_2674_symbol <= Xexit_2676_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_568/simple_obj_ref_565_complete
        Xexit_2670_symbol <= assign_stmt_568_completed_x_x2672_symbol; -- transition branch_block_stmt_513/assign_stmt_568/$exit
        assign_stmt_568_2668_symbol <= Xexit_2670_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_568
      assign_stmt_572_to_assign_stmt_581_2679: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581 
        signal assign_stmt_572_to_assign_stmt_581_2679_start: Boolean;
        signal Xentry_2680_symbol: Boolean;
        signal Xexit_2681_symbol: Boolean;
        signal assign_stmt_572_active_x_x2682_symbol : Boolean;
        signal assign_stmt_572_completed_x_x2683_symbol : Boolean;
        signal ptr_deref_571_trigger_x_x2684_symbol : Boolean;
        signal ptr_deref_571_active_x_x2685_symbol : Boolean;
        signal ptr_deref_571_base_address_calculated_2686_symbol : Boolean;
        signal ptr_deref_571_root_address_calculated_2687_symbol : Boolean;
        signal ptr_deref_571_word_address_calculated_2688_symbol : Boolean;
        signal ptr_deref_571_request_2689_symbol : Boolean;
        signal ptr_deref_571_complete_2700_symbol : Boolean;
        signal assign_stmt_576_active_x_x2713_symbol : Boolean;
        signal assign_stmt_576_completed_x_x2714_symbol : Boolean;
        signal type_cast_575_active_x_x2715_symbol : Boolean;
        signal type_cast_575_trigger_x_x2716_symbol : Boolean;
        signal simple_obj_ref_574_complete_2717_symbol : Boolean;
        signal type_cast_575_complete_2718_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_572_to_assign_stmt_581_2679_start <= assign_stmt_572_to_assign_stmt_581_x_xentry_x_xx_x2468_symbol; -- control passed to block
        Xentry_2680_symbol  <= assign_stmt_572_to_assign_stmt_581_2679_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/$entry
        assign_stmt_572_active_x_x2682_symbol <= ptr_deref_571_complete_2700_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_572_active_
        assign_stmt_572_completed_x_x2683_symbol <= assign_stmt_572_active_x_x2682_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_572_completed_
        ptr_deref_571_trigger_x_x2684_symbol <= ptr_deref_571_word_address_calculated_2688_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_trigger_
        ptr_deref_571_active_x_x2685_symbol <= ptr_deref_571_request_2689_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_active_
        ptr_deref_571_base_address_calculated_2686_symbol <= Xentry_2680_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_base_address_calculated
        ptr_deref_571_root_address_calculated_2687_symbol <= Xentry_2680_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_root_address_calculated
        ptr_deref_571_word_address_calculated_2688_symbol <= ptr_deref_571_root_address_calculated_2687_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_word_address_calculated
        ptr_deref_571_request_2689: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request 
          signal ptr_deref_571_request_2689_start: Boolean;
          signal Xentry_2690_symbol: Boolean;
          signal Xexit_2691_symbol: Boolean;
          signal word_access_2692_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_571_request_2689_start <= ptr_deref_571_trigger_x_x2684_symbol; -- control passed to block
          Xentry_2690_symbol  <= ptr_deref_571_request_2689_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/$entry
          word_access_2692: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access 
            signal word_access_2692_start: Boolean;
            signal Xentry_2693_symbol: Boolean;
            signal Xexit_2694_symbol: Boolean;
            signal word_access_0_2695_symbol : Boolean;
            -- 
          begin -- 
            word_access_2692_start <= Xentry_2690_symbol; -- control passed to block
            Xentry_2693_symbol  <= word_access_2692_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/$entry
            word_access_0_2695: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0 
              signal word_access_0_2695_start: Boolean;
              signal Xentry_2696_symbol: Boolean;
              signal Xexit_2697_symbol: Boolean;
              signal rr_2698_symbol : Boolean;
              signal ra_2699_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2695_start <= Xentry_2693_symbol; -- control passed to block
              Xentry_2696_symbol  <= word_access_0_2695_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/$entry
              rr_2698_symbol <= Xentry_2696_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/rr
              ptr_deref_571_load_0_req_0 <= rr_2698_symbol; -- link to DP
              ra_2699_symbol <= ptr_deref_571_load_0_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/ra
              Xexit_2697_symbol <= ra_2699_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0/$exit
              word_access_0_2695_symbol <= Xexit_2697_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/word_access_0
            Xexit_2694_symbol <= word_access_0_2695_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access/$exit
            word_access_2692_symbol <= Xexit_2694_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/word_access
          Xexit_2691_symbol <= word_access_2692_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request/$exit
          ptr_deref_571_request_2689_symbol <= Xexit_2691_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_request
        ptr_deref_571_complete_2700: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete 
          signal ptr_deref_571_complete_2700_start: Boolean;
          signal Xentry_2701_symbol: Boolean;
          signal Xexit_2702_symbol: Boolean;
          signal word_access_2703_symbol : Boolean;
          signal merge_req_2711_symbol : Boolean;
          signal merge_ack_2712_symbol : Boolean;
          -- 
        begin -- 
          ptr_deref_571_complete_2700_start <= ptr_deref_571_active_x_x2685_symbol; -- control passed to block
          Xentry_2701_symbol  <= ptr_deref_571_complete_2700_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/$entry
          word_access_2703: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access 
            signal word_access_2703_start: Boolean;
            signal Xentry_2704_symbol: Boolean;
            signal Xexit_2705_symbol: Boolean;
            signal word_access_0_2706_symbol : Boolean;
            -- 
          begin -- 
            word_access_2703_start <= Xentry_2701_symbol; -- control passed to block
            Xentry_2704_symbol  <= word_access_2703_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/$entry
            word_access_0_2706: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0 
              signal word_access_0_2706_start: Boolean;
              signal Xentry_2707_symbol: Boolean;
              signal Xexit_2708_symbol: Boolean;
              signal cr_2709_symbol : Boolean;
              signal ca_2710_symbol : Boolean;
              -- 
            begin -- 
              word_access_0_2706_start <= Xentry_2704_symbol; -- control passed to block
              Xentry_2707_symbol  <= word_access_0_2706_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/$entry
              cr_2709_symbol <= Xentry_2707_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/cr
              ptr_deref_571_load_0_req_1 <= cr_2709_symbol; -- link to DP
              ca_2710_symbol <= ptr_deref_571_load_0_ack_1; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/ca
              Xexit_2708_symbol <= ca_2710_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0/$exit
              word_access_0_2706_symbol <= Xexit_2708_symbol; -- control passed from block 
              -- 
            end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/word_access_0
            Xexit_2705_symbol <= word_access_0_2706_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access/$exit
            word_access_2703_symbol <= Xexit_2705_symbol; -- control passed from block 
            -- 
          end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/word_access
          merge_req_2711_symbol <= word_access_2703_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/merge_req
          ptr_deref_571_gather_scatter_req_0 <= merge_req_2711_symbol; -- link to DP
          merge_ack_2712_symbol <= ptr_deref_571_gather_scatter_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/merge_ack
          Xexit_2702_symbol <= merge_ack_2712_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete/$exit
          ptr_deref_571_complete_2700_symbol <= Xexit_2702_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/ptr_deref_571_complete
        assign_stmt_576_active_x_x2713_symbol <= type_cast_575_complete_2718_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_576_active_
        assign_stmt_576_completed_x_x2714_symbol <= assign_stmt_576_active_x_x2713_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/assign_stmt_576_completed_
        type_cast_575_active_x_x2715_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_active_ 
          signal type_cast_575_active_x_x2715_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_575_active_x_x2715_predecessors(0) <= type_cast_575_trigger_x_x2716_symbol;
          type_cast_575_active_x_x2715_predecessors(1) <= simple_obj_ref_574_complete_2717_symbol;
          type_cast_575_active_x_x2715_join: join -- 
            port map( -- 
              preds => type_cast_575_active_x_x2715_predecessors,
              symbol_out => type_cast_575_active_x_x2715_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_active_
        type_cast_575_trigger_x_x2716_symbol <= Xentry_2680_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_trigger_
        simple_obj_ref_574_complete_2717_symbol <= assign_stmt_572_completed_x_x2683_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/simple_obj_ref_574_complete
        type_cast_575_complete_2718: Block -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete 
          signal type_cast_575_complete_2718_start: Boolean;
          signal Xentry_2719_symbol: Boolean;
          signal Xexit_2720_symbol: Boolean;
          signal req_2721_symbol : Boolean;
          signal ack_2722_symbol : Boolean;
          -- 
        begin -- 
          type_cast_575_complete_2718_start <= type_cast_575_active_x_x2715_symbol; -- control passed to block
          Xentry_2719_symbol  <= type_cast_575_complete_2718_start; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/$entry
          req_2721_symbol <= Xentry_2719_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/req
          type_cast_575_inst_req_0 <= req_2721_symbol; -- link to DP
          ack_2722_symbol <= type_cast_575_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/ack
          Xexit_2720_symbol <= ack_2722_symbol; -- transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete/$exit
          type_cast_575_complete_2718_symbol <= Xexit_2720_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/type_cast_575_complete
        Xexit_2681_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/$exit 
          signal Xexit_2681_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          Xexit_2681_predecessors(0) <= ptr_deref_571_base_address_calculated_2686_symbol;
          Xexit_2681_predecessors(1) <= assign_stmt_576_completed_x_x2714_symbol;
          Xexit_2681_join: join -- 
            port map( -- 
              preds => Xexit_2681_predecessors,
              symbol_out => Xexit_2681_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581/$exit
        assign_stmt_572_to_assign_stmt_581_2679_symbol <= Xexit_2681_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_572_to_assign_stmt_581
      assign_stmt_585_2723: Block -- branch_block_stmt_513/assign_stmt_585 
        signal assign_stmt_585_2723_start: Boolean;
        signal Xentry_2724_symbol: Boolean;
        signal Xexit_2725_symbol: Boolean;
        signal assign_stmt_585_active_x_x2726_symbol : Boolean;
        signal assign_stmt_585_completed_x_x2727_symbol : Boolean;
        signal type_cast_584_active_x_x2728_symbol : Boolean;
        signal type_cast_584_trigger_x_x2729_symbol : Boolean;
        signal simple_obj_ref_583_complete_2730_symbol : Boolean;
        signal type_cast_584_complete_2731_symbol : Boolean;
        signal simple_obj_ref_582_trigger_x_x2736_symbol : Boolean;
        signal simple_obj_ref_582_complete_2737_symbol : Boolean;
        -- 
      begin -- 
        assign_stmt_585_2723_start <= assign_stmt_585_x_xentry_x_xx_x2470_symbol; -- control passed to block
        Xentry_2724_symbol  <= assign_stmt_585_2723_start; -- transition branch_block_stmt_513/assign_stmt_585/$entry
        assign_stmt_585_active_x_x2726_symbol <= type_cast_584_complete_2731_symbol; -- transition branch_block_stmt_513/assign_stmt_585/assign_stmt_585_active_
        assign_stmt_585_completed_x_x2727_symbol <= simple_obj_ref_582_complete_2737_symbol; -- transition branch_block_stmt_513/assign_stmt_585/assign_stmt_585_completed_
        type_cast_584_active_x_x2728_block : Block -- non-trivial join transition branch_block_stmt_513/assign_stmt_585/type_cast_584_active_ 
          signal type_cast_584_active_x_x2728_predecessors: BooleanArray(1 downto 0);
          -- 
        begin -- 
          type_cast_584_active_x_x2728_predecessors(0) <= type_cast_584_trigger_x_x2729_symbol;
          type_cast_584_active_x_x2728_predecessors(1) <= simple_obj_ref_583_complete_2730_symbol;
          type_cast_584_active_x_x2728_join: join -- 
            port map( -- 
              preds => type_cast_584_active_x_x2728_predecessors,
              symbol_out => type_cast_584_active_x_x2728_symbol,
              clk => clk,
              reset => reset); -- 
          -- 
        end Block; -- non-trivial join transition branch_block_stmt_513/assign_stmt_585/type_cast_584_active_
        type_cast_584_trigger_x_x2729_symbol <= Xentry_2724_symbol; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_trigger_
        simple_obj_ref_583_complete_2730_symbol <= Xentry_2724_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_583_complete
        type_cast_584_complete_2731: Block -- branch_block_stmt_513/assign_stmt_585/type_cast_584_complete 
          signal type_cast_584_complete_2731_start: Boolean;
          signal Xentry_2732_symbol: Boolean;
          signal Xexit_2733_symbol: Boolean;
          signal req_2734_symbol : Boolean;
          signal ack_2735_symbol : Boolean;
          -- 
        begin -- 
          type_cast_584_complete_2731_start <= type_cast_584_active_x_x2728_symbol; -- control passed to block
          Xentry_2732_symbol  <= type_cast_584_complete_2731_start; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/$entry
          req_2734_symbol <= Xentry_2732_symbol; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/req
          type_cast_584_inst_req_0 <= req_2734_symbol; -- link to DP
          ack_2735_symbol <= type_cast_584_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/ack
          Xexit_2733_symbol <= ack_2735_symbol; -- transition branch_block_stmt_513/assign_stmt_585/type_cast_584_complete/$exit
          type_cast_584_complete_2731_symbol <= Xexit_2733_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_585/type_cast_584_complete
        simple_obj_ref_582_trigger_x_x2736_symbol <= assign_stmt_585_active_x_x2726_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_trigger_
        simple_obj_ref_582_complete_2737: Block -- branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete 
          signal simple_obj_ref_582_complete_2737_start: Boolean;
          signal Xentry_2738_symbol: Boolean;
          signal Xexit_2739_symbol: Boolean;
          signal pipe_wreq_2740_symbol : Boolean;
          signal pipe_wack_2741_symbol : Boolean;
          -- 
        begin -- 
          simple_obj_ref_582_complete_2737_start <= simple_obj_ref_582_trigger_x_x2736_symbol; -- control passed to block
          Xentry_2738_symbol  <= simple_obj_ref_582_complete_2737_start; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/$entry
          pipe_wreq_2740_symbol <= Xentry_2738_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/pipe_wreq
          simple_obj_ref_582_inst_req_0 <= pipe_wreq_2740_symbol; -- link to DP
          pipe_wack_2741_symbol <= simple_obj_ref_582_inst_ack_0; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/pipe_wack
          Xexit_2739_symbol <= pipe_wack_2741_symbol; -- transition branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete/$exit
          simple_obj_ref_582_complete_2737_symbol <= Xexit_2739_symbol; -- control passed from block 
          -- 
        end Block; -- branch_block_stmt_513/assign_stmt_585/simple_obj_ref_582_complete
        Xexit_2725_symbol <= assign_stmt_585_completed_x_x2727_symbol; -- transition branch_block_stmt_513/assign_stmt_585/$exit
        assign_stmt_585_2723_symbol <= Xexit_2725_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/assign_stmt_585
      bb_0_bb_1_PhiReq_2742: Block -- branch_block_stmt_513/bb_0_bb_1_PhiReq 
        signal bb_0_bb_1_PhiReq_2742_start: Boolean;
        signal Xentry_2743_symbol: Boolean;
        signal Xexit_2744_symbol: Boolean;
        -- 
      begin -- 
        bb_0_bb_1_PhiReq_2742_start <= bb_0_bb_1_2454_symbol; -- control passed to block
        Xentry_2743_symbol  <= bb_0_bb_1_PhiReq_2742_start; -- transition branch_block_stmt_513/bb_0_bb_1_PhiReq/$entry
        Xexit_2744_symbol <= Xentry_2743_symbol; -- transition branch_block_stmt_513/bb_0_bb_1_PhiReq/$exit
        bb_0_bb_1_PhiReq_2742_symbol <= Xexit_2744_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/bb_0_bb_1_PhiReq
      bb_1_bb_1_PhiReq_2745: Block -- branch_block_stmt_513/bb_1_bb_1_PhiReq 
        signal bb_1_bb_1_PhiReq_2745_start: Boolean;
        signal Xentry_2746_symbol: Boolean;
        signal Xexit_2747_symbol: Boolean;
        -- 
      begin -- 
        bb_1_bb_1_PhiReq_2745_start <= bb_1_bb_1_2472_symbol; -- control passed to block
        Xentry_2746_symbol  <= bb_1_bb_1_PhiReq_2745_start; -- transition branch_block_stmt_513/bb_1_bb_1_PhiReq/$entry
        Xexit_2747_symbol <= Xentry_2746_symbol; -- transition branch_block_stmt_513/bb_1_bb_1_PhiReq/$exit
        bb_1_bb_1_PhiReq_2745_symbol <= Xexit_2747_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/bb_1_bb_1_PhiReq
      merge_stmt_520_PhiReqMerge_2748_symbol  <=  bb_0_bb_1_PhiReq_2742_symbol or bb_1_bb_1_PhiReq_2745_symbol; -- place branch_block_stmt_513/merge_stmt_520_PhiReqMerge (optimized away) 
      merge_stmt_520_PhiAck_2749: Block -- branch_block_stmt_513/merge_stmt_520_PhiAck 
        signal merge_stmt_520_PhiAck_2749_start: Boolean;
        signal Xentry_2750_symbol: Boolean;
        signal Xexit_2751_symbol: Boolean;
        signal dummy_2752_symbol : Boolean;
        -- 
      begin -- 
        merge_stmt_520_PhiAck_2749_start <= merge_stmt_520_PhiReqMerge_2748_symbol; -- control passed to block
        Xentry_2750_symbol  <= merge_stmt_520_PhiAck_2749_start; -- transition branch_block_stmt_513/merge_stmt_520_PhiAck/$entry
        dummy_2752_symbol <= Xentry_2750_symbol; -- transition branch_block_stmt_513/merge_stmt_520_PhiAck/dummy
        Xexit_2751_symbol <= dummy_2752_symbol; -- transition branch_block_stmt_513/merge_stmt_520_PhiAck/$exit
        merge_stmt_520_PhiAck_2749_symbol <= Xexit_2751_symbol; -- control passed from block 
        -- 
      end Block; -- branch_block_stmt_513/merge_stmt_520_PhiAck
      Xexit_2449_symbol <= branch_block_stmt_513_x_xexit_x_xx_x2451_symbol; -- transition branch_block_stmt_513/$exit
      branch_block_stmt_513_2447_symbol <= Xexit_2449_symbol; -- control passed from block 
      -- 
    end Block; -- branch_block_stmt_513
    Xexit_2446_symbol <= branch_block_stmt_513_2447_symbol; -- transition $exit
    fin  <=  '1' when Xexit_2446_symbol else '0'; -- fin symbol when control-path exits
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_545_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_545_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_545_root_address : std_logic_vector(2 downto 0);
    signal iNsTr_10_564 : std_logic_vector(31 downto 0);
    signal iNsTr_12_572 : std_logic_vector(31 downto 0);
    signal iNsTr_13_576 : std_logic_vector(31 downto 0);
    signal iNsTr_14_581 : std_logic_vector(31 downto 0);
    signal iNsTr_1_525 : std_logic_vector(31 downto 0);
    signal iNsTr_2_529 : std_logic_vector(31 downto 0);
    signal iNsTr_3_533 : std_logic_vector(31 downto 0);
    signal iNsTr_5_541 : std_logic_vector(31 downto 0);
    signal iNsTr_6_546 : std_logic_vector(31 downto 0);
    signal iNsTr_7_550 : std_logic_vector(31 downto 0);
    signal iNsTr_8_555 : std_logic_vector(31 downto 0);
    signal lptr_518 : std_logic_vector(31 downto 0);
    signal ptr_deref_535_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_535_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_535_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_540_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_540_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_549_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_549_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_549_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_549_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_549_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_571_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_571_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_527_wire : std_logic_vector(31 downto 0);
    signal type_cast_558_wire : std_logic_vector(31 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_584_wire : std_logic_vector(31 downto 0);
    signal xxoutput_modulexxbodyxxlptr_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_545_final_offset <= "001";
    iNsTr_10_564 <= "00000000000000000000000000000000";
    iNsTr_14_581 <= "00000000000000000000000000000000";
    iNsTr_1_525 <= "00000000000000000000000000000000";
    iNsTr_8_555 <= "00000000000000000000000000000000";
    lptr_518 <= "00000000000000000000000000000000";
    ptr_deref_535_word_address_0 <= "0";
    ptr_deref_540_word_address_0 <= "0";
    ptr_deref_549_word_offset_0 <= "000";
    ptr_deref_571_word_address_0 <= "0";
    type_cast_567_wire_constant <= "00000001";
    xxoutput_modulexxbodyxxlptr_alloc_base_address <= "0";
    array_obj_ref_545_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_5_541, dout => array_obj_ref_545_resized_base_address, req => array_obj_ref_545_base_resize_req_0, ack => array_obj_ref_545_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_545_final_reg: RegisterBase generic map(in_data_width => 3,out_data_width => 32) -- 
      port map( din => array_obj_ref_545_root_address, dout => iNsTr_6_546, req => array_obj_ref_545_final_reg_req_0, ack => array_obj_ref_545_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_549_base_resize: RegisterBase generic map(in_data_width => 32,out_data_width => 3) -- 
      port map( din => iNsTr_6_546, dout => ptr_deref_549_resized_base_address, req => ptr_deref_549_base_resize_req_0, ack => ptr_deref_549_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_528_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => simple_obj_ref_527_wire, dout => iNsTr_2_529, req => type_cast_528_inst_req_0, ack => type_cast_528_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_532_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_2_529, dout => iNsTr_3_533, req => type_cast_532_inst_req_0, ack => type_cast_532_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_558_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_7_550, dout => type_cast_558_wire, req => type_cast_558_inst_req_0, ack => type_cast_558_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_575_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_12_572, dout => iNsTr_13_576, req => type_cast_575_inst_req_0, ack => type_cast_575_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_584_inst: RegisterBase generic map(in_data_width => 32,out_data_width => 32) -- 
      port map( din => iNsTr_13_576, dout => type_cast_584_wire, req => type_cast_584_inst_req_0, ack => type_cast_584_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_535_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_535_gather_scatter_ack_0 <= ptr_deref_535_gather_scatter_req_0;
      aggregated_sig <= iNsTr_3_533;
      ptr_deref_535_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_540_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_540_gather_scatter_ack_0 <= ptr_deref_540_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_540_data_0;
      iNsTr_5_541 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_549_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_549_addr_0_ack_0 <= ptr_deref_549_addr_0_req_0;
      aggregated_sig <= ptr_deref_549_root_address;
      ptr_deref_549_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_549_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_549_gather_scatter_ack_0 <= ptr_deref_549_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_549_data_0;
      iNsTr_7_550 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_549_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_549_root_address_inst_ack_0 <= ptr_deref_549_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_549_resized_base_address;
      ptr_deref_549_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_571_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_571_gather_scatter_ack_0 <= ptr_deref_571_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_571_data_0;
      iNsTr_12_572 <= aggregated_sig(31 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_545_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_545_resized_base_address;
      array_obj_ref_545_root_address <= data_out(2 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "001",
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_545_root_address_inst_req_0,
          ackL => array_obj_ref_545_root_address_inst_ack_0,
          reqR => array_obj_ref_545_root_address_inst_req_1,
          ackR => array_obj_ref_545_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared load operator group (0) : ptr_deref_540_load_0 ptr_deref_571_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_540_load_0_req_0;
      reqL(0) <= ptr_deref_571_load_0_req_0;
      ptr_deref_540_load_0_ack_0 <= ackL(1);
      ptr_deref_571_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_540_load_0_req_1;
      reqR(0) <= ptr_deref_571_load_0_req_1;
      ptr_deref_540_load_0_ack_1 <= ackR(1);
      ptr_deref_571_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_540_word_address_0 & ptr_deref_571_word_address_0;
      ptr_deref_540_data_0 <= data_out(63 downto 32);
      ptr_deref_571_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_17_lr_req(0),
          mack => memory_space_17_lr_ack(0),
          maddr => memory_space_17_lr_addr(0 downto 0),
          mtag => memory_space_17_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_17_lc_req(0),
          mack => memory_space_17_lc_ack(0),
          mdata => memory_space_17_lc_data(31 downto 0),
          mtag => memory_space_17_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_549_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_549_load_0_req_0;
      ptr_deref_549_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_549_load_0_req_1;
      ptr_deref_549_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_549_word_address_0;
      ptr_deref_549_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 3,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(2 downto 0),
          mtag => memory_space_1_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_535_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_535_store_0_req_0;
      ptr_deref_535_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_535_store_0_req_1;
      ptr_deref_535_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_535_word_address_0;
      data_in <= ptr_deref_535_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_17_sr_req(0),
          mack => memory_space_17_sr_ack(0),
          maddr => memory_space_17_sr_addr(0 downto 0),
          mdata => memory_space_17_sr_data(31 downto 0),
          mtag => memory_space_17_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_17_sc_req(0),
          mack => memory_space_17_sc_ack(0),
          mtag => memory_space_17_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_527_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_527_inst_req_0;
      simple_obj_ref_527_inst_ack_0 <= ack(0);
      simple_obj_ref_527_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => foo_out_pipe_read_req(0),
          oack => foo_out_pipe_read_ack(0),
          odata => foo_out_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : simple_obj_ref_556_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_556_inst_req_0;
      simple_obj_ref_556_inst_ack_0 <= ack(0);
      data_in <= type_cast_558_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => output_data_pipe_write_req(0),
          oack => output_data_pipe_write_ack(0),
          odata => output_data_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_565_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_565_inst_req_0;
      simple_obj_ref_565_inst_ack_0 <= ack(0);
      data_in <= type_cast_567_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_582_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_582_inst_req_0;
      simple_obj_ref_582_inst_ack_0 <= ack(0);
      data_in <= type_cast_584_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_put_pipe_write_req(0),
          oack => free_queue_put_pipe_write_ack(0),
          odata => free_queue_put_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  RegisterBank_memory_space_17: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_17_lr_addr,
      lr_req_in => memory_space_17_lr_req,
      lr_ack_out => memory_space_17_lr_ack,
      lr_tag_in => memory_space_17_lr_tag,
      lc_req_in => memory_space_17_lc_req,
      lc_ack_out => memory_space_17_lc_ack,
      lc_data_out => memory_space_17_lc_data,
      lc_tag_out => memory_space_17_lc_tag,
      sr_addr_in => memory_space_17_sr_addr,
      sr_data_in => memory_space_17_sr_data,
      sr_req_in => memory_space_17_sr_req,
      sr_ack_out => memory_space_17_sr_ack,
      sr_tag_in => memory_space_17_sr_tag,
      sc_req_in=> memory_space_17_sc_req,
      sc_ack_out => memory_space_17_sc_ack,
      sc_tag_out => memory_space_17_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity test_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    input_data_pipe_write_data: in std_logic_vector(31 downto 0);
    input_data_pipe_write_req : in std_logic_vector(0 downto 0);
    input_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    output_data_pipe_read_data: out std_logic_vector(31 downto 0);
    output_data_pipe_read_req : in std_logic_vector(0 downto 0);
    output_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of test_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(2 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(2 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(2 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(95 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(2 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(95 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(2 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(2 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(5 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(1 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  -- interface signals to connect to memory space memory_space_4
  -- interface signals to connect to memory space memory_space_5
  -- interface signals to connect to memory space memory_space_6
  -- interface signals to connect to memory space memory_space_7
  -- interface signals to connect to memory space memory_space_8
  -- interface signals to connect to memory space memory_space_9
  -- declarations related to module foo
  component foo is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      foo_in_pipe_read_req : out  std_logic_vector(0 downto 0);
      foo_in_pipe_read_ack : in   std_logic_vector(0 downto 0);
      foo_in_pipe_read_data : in   std_logic_vector(31 downto 0);
      foo_out_pipe_write_req : out  std_logic_vector(0 downto 0);
      foo_out_pipe_write_ack : in   std_logic_vector(0 downto 0);
      foo_out_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module foo
  signal foo_tag_in    : std_logic_vector(0 downto 0);
  signal foo_tag_out   : std_logic_vector(0 downto 0);
  signal foo_start : std_logic;
  signal foo_fin   : std_logic;
  -- declarations related to module free_queue_manager
  component free_queue_manager is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(1 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(1 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(1 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(1 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(1 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module free_queue_manager
  signal free_queue_manager_tag_in    : std_logic_vector(0 downto 0);
  signal free_queue_manager_tag_out   : std_logic_vector(0 downto 0);
  signal free_queue_manager_start : std_logic;
  signal free_queue_manager_fin   : std_logic;
  -- declarations related to module input_module
  component input_module is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(2 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_data_pipe_read_data : in   std_logic_vector(31 downto 0);
      foo_in_pipe_write_req : out  std_logic_vector(0 downto 0);
      foo_in_pipe_write_ack : in   std_logic_vector(0 downto 0);
      foo_in_pipe_write_data : out  std_logic_vector(31 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module input_module
  signal input_module_tag_in    : std_logic_vector(0 downto 0);
  signal input_module_tag_out   : std_logic_vector(0 downto 0);
  signal input_module_start : std_logic;
  signal input_module_fin   : std_logic;
  -- declarations related to module mem_load_x_x
  component mem_load_x_x is -- 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(7 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module mem_load_x_x
  signal mem_load_x_x_address :  std_logic_vector(31 downto 0);
  signal mem_load_x_x_data :  std_logic_vector(7 downto 0);
  signal mem_load_x_x_in_args    : std_logic_vector(31 downto 0);
  signal mem_load_x_x_out_args   : std_logic_vector(7 downto 0);
  signal mem_load_x_x_tag_in    : std_logic_vector(0 downto 0);
  signal mem_load_x_x_tag_out   : std_logic_vector(0 downto 0);
  signal mem_load_x_x_start : std_logic;
  signal mem_load_x_x_fin   : std_logic;
  -- declarations related to module mem_store_x_x
  component mem_store_x_x is -- 
    port ( -- 
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(7 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module mem_store_x_x
  signal mem_store_x_x_address :  std_logic_vector(31 downto 0);
  signal mem_store_x_x_data :  std_logic_vector(7 downto 0);
  signal mem_store_x_x_in_args    : std_logic_vector(39 downto 0);
  signal mem_store_x_x_tag_in    : std_logic_vector(0 downto 0);
  signal mem_store_x_x_tag_out   : std_logic_vector(0 downto 0);
  signal mem_store_x_x_start : std_logic;
  signal mem_store_x_x_fin   : std_logic;
  -- declarations related to module output_module
  component output_module is -- 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      foo_out_pipe_read_req : out  std_logic_vector(0 downto 0);
      foo_out_pipe_read_ack : in   std_logic_vector(0 downto 0);
      foo_out_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      output_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_data_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- argument signals for module output_module
  signal output_module_tag_in    : std_logic_vector(0 downto 0);
  signal output_module_tag_out   : std_logic_vector(0 downto 0);
  signal output_module_start : std_logic;
  signal output_module_fin   : std_logic;
  -- aggregate signals for write to pipe foo_in
  signal foo_in_pipe_write_data: std_logic_vector(31 downto 0);
  signal foo_in_pipe_write_req: std_logic_vector(0 downto 0);
  signal foo_in_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe foo_in
  signal foo_in_pipe_read_data: std_logic_vector(31 downto 0);
  signal foo_in_pipe_read_req: std_logic_vector(0 downto 0);
  signal foo_in_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe foo_out
  signal foo_out_pipe_write_data: std_logic_vector(31 downto 0);
  signal foo_out_pipe_write_req: std_logic_vector(0 downto 0);
  signal foo_out_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe foo_out
  signal foo_out_pipe_read_data: std_logic_vector(31 downto 0);
  signal foo_out_pipe_read_req: std_logic_vector(0 downto 0);
  signal foo_out_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_get
  signal free_queue_get_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_get
  signal free_queue_get_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_put
  signal free_queue_put_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_put
  signal free_queue_put_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_request
  signal free_queue_request_pipe_write_data: std_logic_vector(15 downto 0);
  signal free_queue_request_pipe_write_req: std_logic_vector(1 downto 0);
  signal free_queue_request_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe free_queue_request
  signal free_queue_request_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_request_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_request_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_data
  signal input_data_pipe_read_data: std_logic_vector(31 downto 0);
  signal input_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe output_data
  signal output_data_pipe_write_data: std_logic_vector(31 downto 0);
  signal output_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal output_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module foo
  foo_instance:foo-- 
    port map(-- 
      start => foo_start,
      fin => foo_fin,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(8 downto 6),
      memory_space_1_lr_tag => memory_space_1_lr_tag(5 downto 4),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 4),
      memory_space_1_sr_req => memory_space_1_sr_req(2 downto 2),
      memory_space_1_sr_ack => memory_space_1_sr_ack(2 downto 2),
      memory_space_1_sr_addr => memory_space_1_sr_addr(8 downto 6),
      memory_space_1_sr_data => memory_space_1_sr_data(95 downto 64),
      memory_space_1_sr_tag => memory_space_1_sr_tag(5 downto 4),
      memory_space_1_sc_req => memory_space_1_sc_req(2 downto 2),
      memory_space_1_sc_ack => memory_space_1_sc_ack(2 downto 2),
      memory_space_1_sc_tag => memory_space_1_sc_tag(5 downto 4),
      foo_in_pipe_read_req => foo_in_pipe_read_req(0 downto 0),
      foo_in_pipe_read_ack => foo_in_pipe_read_ack(0 downto 0),
      foo_in_pipe_read_data => foo_in_pipe_read_data(31 downto 0),
      foo_out_pipe_write_req => foo_out_pipe_write_req(0 downto 0),
      foo_out_pipe_write_ack => foo_out_pipe_write_ack(0 downto 0),
      foo_out_pipe_write_data => foo_out_pipe_write_data(31 downto 0),
      tag_in => foo_tag_in,
      tag_out => foo_tag_out-- 
    ); -- 
  -- module will be run forever 
  foo_tag_in <= (others => '0');
  foo_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => foo_start, fin => foo_fin);
  -- module free_queue_manager
  free_queue_manager_instance:free_queue_manager-- 
    port map(-- 
      start => free_queue_manager_start,
      fin => free_queue_manager_fin,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(2 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(1 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(1 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(3 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(1 downto 1),
      memory_space_1_sr_ack => memory_space_1_sr_ack(1 downto 1),
      memory_space_1_sr_addr => memory_space_1_sr_addr(5 downto 3),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 32),
      memory_space_1_sr_tag => memory_space_1_sr_tag(3 downto 2),
      memory_space_1_sc_req => memory_space_1_sc_req(1 downto 1),
      memory_space_1_sc_ack => memory_space_1_sc_ack(1 downto 1),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 2),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(1 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      free_queue_put_pipe_read_req => free_queue_put_pipe_read_req(0 downto 0),
      free_queue_put_pipe_read_ack => free_queue_put_pipe_read_ack(0 downto 0),
      free_queue_put_pipe_read_data => free_queue_put_pipe_read_data(31 downto 0),
      free_queue_request_pipe_read_req => free_queue_request_pipe_read_req(0 downto 0),
      free_queue_request_pipe_read_ack => free_queue_request_pipe_read_ack(0 downto 0),
      free_queue_request_pipe_read_data => free_queue_request_pipe_read_data(7 downto 0),
      free_queue_get_pipe_write_req => free_queue_get_pipe_write_req(0 downto 0),
      free_queue_get_pipe_write_ack => free_queue_get_pipe_write_ack(0 downto 0),
      free_queue_get_pipe_write_data => free_queue_get_pipe_write_data(31 downto 0),
      tag_in => free_queue_manager_tag_in,
      tag_out => free_queue_manager_tag_out-- 
    ); -- 
  -- module will be run forever 
  free_queue_manager_tag_in <= (others => '0');
  free_queue_manager_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => free_queue_manager_start, fin => free_queue_manager_fin);
  -- module input_module
  input_module_instance:input_module-- 
    port map(-- 
      start => input_module_start,
      fin => input_module_fin,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(2 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(1 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      free_queue_get_pipe_read_req => free_queue_get_pipe_read_req(0 downto 0),
      free_queue_get_pipe_read_ack => free_queue_get_pipe_read_ack(0 downto 0),
      free_queue_get_pipe_read_data => free_queue_get_pipe_read_data(31 downto 0),
      input_data_pipe_read_req => input_data_pipe_read_req(0 downto 0),
      input_data_pipe_read_ack => input_data_pipe_read_ack(0 downto 0),
      input_data_pipe_read_data => input_data_pipe_read_data(31 downto 0),
      foo_in_pipe_write_req => foo_in_pipe_write_req(0 downto 0),
      foo_in_pipe_write_ack => foo_in_pipe_write_ack(0 downto 0),
      foo_in_pipe_write_data => foo_in_pipe_write_data(31 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(0 downto 0),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(0 downto 0),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(7 downto 0),
      tag_in => input_module_tag_in,
      tag_out => input_module_tag_out-- 
    ); -- 
  -- module will be run forever 
  input_module_tag_in <= (others => '0');
  input_module_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => input_module_start, fin => input_module_fin);
  -- module mem_load_x_x
  mem_load_x_x_start <= '0';
  mem_load_x_x_instance:mem_load_x_x-- 
    port map(-- 
      address => mem_load_x_x_address,
      data => mem_load_x_x_data,
      start => mem_load_x_x_start,
      fin => mem_load_x_x_fin,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(7 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => mem_load_x_x_tag_in,
      tag_out => mem_load_x_x_tag_out-- 
    ); -- 
  -- module mem_store_x_x
  mem_store_x_x_start <= '0';
  mem_store_x_x_instance:mem_store_x_x-- 
    port map(-- 
      address => mem_store_x_x_address,
      data => mem_store_x_x_data,
      start => mem_store_x_x_start,
      fin => mem_store_x_x_fin,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(0 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(7 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(0 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      tag_in => mem_store_x_x_tag_in,
      tag_out => mem_store_x_x_tag_out-- 
    ); -- 
  -- module output_module
  output_module_instance:output_module-- 
    port map(-- 
      start => output_module_start,
      fin => output_module_fin,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(5 downto 3),
      memory_space_1_lr_tag => memory_space_1_lr_tag(3 downto 2),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 2),
      foo_out_pipe_read_req => foo_out_pipe_read_req(0 downto 0),
      foo_out_pipe_read_ack => foo_out_pipe_read_ack(0 downto 0),
      foo_out_pipe_read_data => foo_out_pipe_read_data(31 downto 0),
      free_queue_put_pipe_write_req => free_queue_put_pipe_write_req(0 downto 0),
      free_queue_put_pipe_write_ack => free_queue_put_pipe_write_ack(0 downto 0),
      free_queue_put_pipe_write_data => free_queue_put_pipe_write_data(31 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(1 downto 1),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(1 downto 1),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(15 downto 8),
      output_data_pipe_write_req => output_data_pipe_write_req(0 downto 0),
      output_data_pipe_write_ack => output_data_pipe_write_ack(0 downto 0),
      output_data_pipe_write_data => output_data_pipe_write_data(31 downto 0),
      tag_in => output_module_tag_in,
      tag_out => output_module_tag_out-- 
    ); -- 
  -- module will be run forever 
  output_module_tag_in <= (others => '0');
  output_module_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start => output_module_start, fin => output_module_fin);
  foo_in_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => foo_in_pipe_read_req,
      read_ack => foo_in_pipe_read_ack,
      read_data => foo_in_pipe_read_data,
      write_req => foo_in_pipe_write_req,
      write_ack => foo_in_pipe_write_ack,
      write_data => foo_in_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  foo_out_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => foo_out_pipe_read_req,
      read_ack => foo_out_pipe_read_ack,
      read_data => foo_out_pipe_read_data,
      write_req => foo_out_pipe_write_req,
      write_ack => foo_out_pipe_write_ack,
      write_data => foo_out_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_get_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_get_pipe_read_req,
      read_ack => free_queue_get_pipe_read_ack,
      read_data => free_queue_get_pipe_read_data,
      write_req => free_queue_get_pipe_write_req,
      write_ack => free_queue_get_pipe_write_ack,
      write_data => free_queue_get_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_put_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_put_pipe_read_req,
      read_ack => free_queue_put_pipe_read_ack,
      read_data => free_queue_put_pipe_read_data,
      write_req => free_queue_put_pipe_write_req,
      write_ack => free_queue_put_pipe_write_ack,
      write_data => free_queue_put_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_request_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_request_pipe_read_req,
      read_ack => free_queue_request_pipe_read_ack,
      read_data => free_queue_request_pipe_read_data,
      write_req => free_queue_request_pipe_write_req,
      write_ack => free_queue_request_pipe_write_ack,
      write_data => free_queue_request_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => input_data_pipe_read_req,
      read_ack => input_data_pipe_read_ack,
      read_data => input_data_pipe_read_data,
      write_req => input_data_pipe_write_req,
      write_ack => input_data_pipe_write_ack,
      write_data => input_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  output_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => output_data_pipe_read_req,
      read_ack => output_data_pipe_read_ack,
      read_data => output_data_pipe_read_data,
      write_req => output_data_pipe_write_req,
      write_ack => output_data_pipe_write_ack,
      write_data => output_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  RegisterBank_memory_space_0: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 1,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_1: register_bank -- 
    generic map(-- 
      num_loads => 3,
      num_stores => 3,
      addr_width => 3,
      data_width => 32,
      tag_width => 2,
      num_registers => 4) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_2: register_bank -- 
    generic map(-- 
      num_loads => 2,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      num_registers => 1) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
use work.Utility_Package.all;
use work.Vhpi_Foreign.all;
entity test_system_Test_Bench is -- 
  -- 
end entity;
architecture VhpiLink of test_system_Test_Bench is -- 
  component test_system is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      input_data_pipe_write_data: in std_logic_vector(31 downto 0);
      input_data_pipe_write_req : in std_logic_vector(0 downto 0);
      input_data_pipe_write_ack : out std_logic_vector(0 downto 0);
      output_data_pipe_read_data: out std_logic_vector(31 downto 0);
      output_data_pipe_read_req : in std_logic_vector(0 downto 0);
      output_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
    -- 
  end component;
  signal clk: std_logic := '0';
  signal reset: std_logic := '1';
  signal foo_tag_in: std_logic_vector(0 downto 0);
  signal foo_tag_out: std_logic_vector(0 downto 0);
  signal foo_start : std_logic := '0';
  signal foo_fin   : std_logic := '0';
  signal free_queue_manager_tag_in: std_logic_vector(0 downto 0);
  signal free_queue_manager_tag_out: std_logic_vector(0 downto 0);
  signal free_queue_manager_start : std_logic := '0';
  signal free_queue_manager_fin   : std_logic := '0';
  signal input_module_tag_in: std_logic_vector(0 downto 0);
  signal input_module_tag_out: std_logic_vector(0 downto 0);
  signal input_module_start : std_logic := '0';
  signal input_module_fin   : std_logic := '0';
  signal output_module_tag_in: std_logic_vector(0 downto 0);
  signal output_module_tag_out: std_logic_vector(0 downto 0);
  signal output_module_start : std_logic := '0';
  signal output_module_fin   : std_logic := '0';
  -- write to pipe input_data
  signal input_data_pipe_write_data: std_logic_vector(31 downto 0);
  signal input_data_pipe_write_req : std_logic_vector(0 downto 0) := (others => '0');
  signal input_data_pipe_write_ack : std_logic_vector(0 downto 0);
  -- read from pipe output_data
  signal output_data_pipe_read_data: std_logic_vector(31 downto 0);
  signal output_data_pipe_read_req : std_logic_vector(0 downto 0) := (others => '0');
  signal output_data_pipe_read_ack : std_logic_vector(0 downto 0);
  -- 
begin --
  -- clock/reset generation 
  clk <= not clk after 5 ns;
  process
  begin --
    Vhpi_Initialize;
    wait until clk = '1';
    reset <= '0';
    while true loop --
      wait until clk = '0';
      Vhpi_Listen;
      Vhpi_Send;
      --
    end loop;
    wait;
    --
  end process;
  -- connect all the top-level modules to Vhpi
  process
  variable val_string, obj_ref: VhpiString;
  begin --
    wait until reset = '0';
    while true loop -- 
      wait until clk = '0';
      wait for 1 ns; 
      obj_ref := Pack_String_To_Vhpi_String("input_data req");
      Vhpi_Get_Port_Value(obj_ref,val_string,1);
      input_data_pipe_write_req <= Unpack_String(val_string,1);
      obj_ref := Pack_String_To_Vhpi_String("input_data 0");
      Vhpi_Get_Port_Value(obj_ref,val_string,32);
      input_data_pipe_write_data <= Unpack_String(val_string,32);
      wait until clk = '1';
      obj_ref := Pack_String_To_Vhpi_String("input_data ack");
      val_string := Pack_SLV_To_Vhpi_String(input_data_pipe_write_ack);
      Vhpi_Set_Port_Value(obj_ref,val_string,1);
      -- 
    end loop;
    --
  end process;
  process
  variable val_string, obj_ref: VhpiString;
  begin --
    wait until reset = '0';
    while true loop -- 
      wait until clk = '0';
      wait for 1 ns; 
      obj_ref := Pack_String_To_Vhpi_String("output_data req");
      Vhpi_Get_Port_Value(obj_ref,val_string,1);
      output_data_pipe_read_req <= Unpack_String(val_string,1);
      wait until clk = '1';
      obj_ref := Pack_String_To_Vhpi_String("output_data ack");
      val_string := Pack_SLV_To_Vhpi_String(output_data_pipe_read_ack);
      Vhpi_Set_Port_Value(obj_ref,val_string,1);
      obj_ref := Pack_String_To_Vhpi_String("output_data 0");
      val_string := Pack_SLV_To_Vhpi_String(output_data_pipe_read_data);
      Vhpi_Set_Port_Value(obj_ref,val_string,32);
      -- 
    end loop;
    --
  end process;
  test_system_instance: test_system -- 
    port map ( -- 
      clk => clk,
      reset => reset,
      input_data_pipe_write_data  => input_data_pipe_write_data, 
      input_data_pipe_write_req  => input_data_pipe_write_req, 
      input_data_pipe_write_ack  => input_data_pipe_write_ack,
      output_data_pipe_read_data  => output_data_pipe_read_data, 
      output_data_pipe_read_req  => output_data_pipe_read_req, 
      output_data_pipe_read_ack  => output_data_pipe_read_ack ); -- 
  -- 
end VhpiLink;
